----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 5/24/2019 11:15:35 AM
-- Design Name: 
-- Module Name: exp_fun - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------



library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity exp_fun is
    Port ( clk : in std_logic;
           inp_wt : in STD_LOGIC_VECTOR (19 downto 0);
           out_wt : out STD_LOGIC_VECTOR (15 downto 0));
end exp_fun;

architecture Behavioral of exp_fun is
signal sig_inp: STD_LOGIC_VECTOR (19 downto 0);
signal sig_out: STD_LOGIC_VECTOR (15 downto 0);
begin

process(clk)
begin
if clk'event and clk = '0' then 
    out_wt <= sig_out;
end if;

end process;

sig_inp <= inp_wt;


----------------------------------------------------------------------------------------------------------------------------------------------------------------
--------------------------------- E.X.P.O.N.E.N.T C.A.L.C.U.L.A.T.I.O.N ----------------------------------------------------------------------------------------
----------------------------------------------------------------------------------------------------------------------------------------------------------------
----------------
--"Sigma_r = 5"
--"a = 3"
-----------------------------
sig_out <= 
"1000000000000000" when sig_inp  = "00000000000000000000" else
"0111111101101110" when sig_inp <= "00000000000000000001" else
"0111111011011110" when sig_inp <= "00000000000000000010" else
"0111111001001101" when sig_inp <= "00000000000000000011" else
"0111110110111110" when sig_inp <= "00000000000000000100" else
"0111110100101111" when sig_inp <= "00000000000000000101" else
"0111110010100001" when sig_inp <= "00000000000000000110" else
"0111110000010100" when sig_inp <= "00000000000000000111" else
"0111101110000111" when sig_inp <= "00000000000000001000" else
"0111101011111011" when sig_inp <= "00000000000000001001" else
"0111101001101111" when sig_inp <= "00000000000000001010" else
"0111100111100100" when sig_inp <= "00000000000000001011" else
"0111100101011010" when sig_inp <= "00000000000000001100" else
"0111100011010000" when sig_inp <= "00000000000000001101" else
"0111100001000111" when sig_inp <= "00000000000000001110" else
"0111011110111110" when sig_inp <= "00000000000000001111" else
"0111011100110110" when sig_inp <= "00000000000000010000" else
"0111011010101111" when sig_inp <= "00000000000000010001" else
"0111011000101000" when sig_inp <= "00000000000000010010" else
"0111010110100010" when sig_inp <= "00000000000000010011" else
"0111010100011100" when sig_inp <= "00000000000000010100" else
"0111010010011000" when sig_inp <= "00000000000000010101" else
"0111010000010011" when sig_inp <= "00000000000000010110" else
"0111001110001111" when sig_inp <= "00000000000000010111" else
"0111001100001100" when sig_inp <= "00000000000000011000" else
"0111001010001010" when sig_inp <= "00000000000000011001" else
"0111001000001000" when sig_inp <= "00000000000000011010" else
"0111000110000110" when sig_inp <= "00000000000000011011" else
"0111000100000101" when sig_inp <= "00000000000000011100" else
"0111000010000101" when sig_inp <= "00000000000000011101" else
"0111000000000101" when sig_inp <= "00000000000000011110" else
"0110111110000110" when sig_inp <= "00000000000000011111" else
"0110111100000111" when sig_inp <= "00000000000000100000" else
"0110111010001001" when sig_inp <= "00000000000000100001" else
"0110111000001100" when sig_inp <= "00000000000000100010" else
"0110110110001111" when sig_inp <= "00000000000000100011" else
"0110110100010011" when sig_inp <= "00000000000000100100" else
"0110110010010111" when sig_inp <= "00000000000000100101" else
"0110110000011011" when sig_inp <= "00000000000000100110" else
"0110101110100001" when sig_inp <= "00000000000000100111" else
"0110101100100111" when sig_inp <= "00000000000000101000" else
"0110101010101101" when sig_inp <= "00000000000000101001" else
"0110101000110100" when sig_inp <= "00000000000000101010" else
"0110100110111011" when sig_inp <= "00000000000000101011" else
"0110100101000011" when sig_inp <= "00000000000000101100" else
"0110100011001100" when sig_inp <= "00000000000000101101" else
"0110100001010101" when sig_inp <= "00000000000000101110" else
"0110011111011110" when sig_inp <= "00000000000000101111" else
"0110011101101000" when sig_inp <= "00000000000000110000" else
"0110011011110011" when sig_inp <= "00000000000000110001" else
"0110011001111110" when sig_inp <= "00000000000000110010" else
"0110011000001010" when sig_inp <= "00000000000000110011" else
"0110010110010110" when sig_inp <= "00000000000000110100" else
"0110010100100011" when sig_inp <= "00000000000000110101" else
"0110010010110000" when sig_inp <= "00000000000000110110" else
"0110010000111101" when sig_inp <= "00000000000000110111" else
"0110001111001100" when sig_inp <= "00000000000000111000" else
"0110001101011010" when sig_inp <= "00000000000000111001" else
"0110001011101010" when sig_inp <= "00000000000000111010" else
"0110001001111001" when sig_inp <= "00000000000000111011" else
"0110001000001001" when sig_inp <= "00000000000000111100" else
"0110000110011010" when sig_inp <= "00000000000000111101" else
"0110000100101011" when sig_inp <= "00000000000000111110" else
"0110000010111101" when sig_inp <= "00000000000000111111" else
"0110000001001111" when sig_inp <= "00000000000001000000" else
"0101111111100010" when sig_inp <= "00000000000001000001" else
"0101111101110101" when sig_inp <= "00000000000001000010" else
"0101111100001001" when sig_inp <= "00000000000001000011" else
"0101111010011101" when sig_inp <= "00000000000001000100" else
"0101111000110001" when sig_inp <= "00000000000001000101" else
"0101110111000110" when sig_inp <= "00000000000001000110" else
"0101110101011100" when sig_inp <= "00000000000001000111" else
"0101110011110010" when sig_inp <= "00000000000001001000" else
"0101110010001000" when sig_inp <= "00000000000001001001" else
"0101110000011111" when sig_inp <= "00000000000001001010" else
"0101101110110111" when sig_inp <= "00000000000001001011" else
"0101101101001111" when sig_inp <= "00000000000001001100" else
"0101101011100111" when sig_inp <= "00000000000001001101" else
"0101101010000000" when sig_inp <= "00000000000001001110" else
"0101101000011001" when sig_inp <= "00000000000001001111" else
"0101100110110011" when sig_inp <= "00000000000001010000" else
"0101100101001101" when sig_inp <= "00000000000001010001" else
"0101100011101000" when sig_inp <= "00000000000001010010" else
"0101100010000011" when sig_inp <= "00000000000001010011" else
"0101100000011110" when sig_inp <= "00000000000001010100" else
"0101011110111010" when sig_inp <= "00000000000001010101" else
"0101011101010111" when sig_inp <= "00000000000001010110" else
"0101011011110011" when sig_inp <= "00000000000001010111" else
"0101011010010001" when sig_inp <= "00000000000001011000" else
"0101011000101110" when sig_inp <= "00000000000001011001" else
"0101010111001101" when sig_inp <= "00000000000001011010" else
"0101010101101011" when sig_inp <= "00000000000001011011" else
"0101010100001010" when sig_inp <= "00000000000001011100" else
"0101010010101010" when sig_inp <= "00000000000001011101" else
"0101010001001010" when sig_inp <= "00000000000001011110" else
"0101001111101010" when sig_inp <= "00000000000001011111" else
"0101001110001011" when sig_inp <= "00000000000001100000" else
"0101001100101100" when sig_inp <= "00000000000001100001" else
"0101001011001101" when sig_inp <= "00000000000001100010" else
"0101001001101111" when sig_inp <= "00000000000001100011" else
"0101001000010010" when sig_inp <= "00000000000001100100" else
"0101000110110101" when sig_inp <= "00000000000001100101" else
"0101000101011000" when sig_inp <= "00000000000001100110" else
"0101000011111011" when sig_inp <= "00000000000001100111" else
"0101000010011111" when sig_inp <= "00000000000001101000" else
"0101000001000100" when sig_inp <= "00000000000001101001" else
"0100111111101001" when sig_inp <= "00000000000001101010" else
"0100111110001110" when sig_inp <= "00000000000001101011" else
"0100111100110100" when sig_inp <= "00000000000001101100" else
"0100111011011010" when sig_inp <= "00000000000001101101" else
"0100111010000000" when sig_inp <= "00000000000001101110" else
"0100111000100111" when sig_inp <= "00000000000001101111" else
"0100110111001111" when sig_inp <= "00000000000001110000" else
"0100110101110110" when sig_inp <= "00000000000001110001" else
"0100110100011110" when sig_inp <= "00000000000001110010" else
"0100110011000111" when sig_inp <= "00000000000001110011" else
"0100110001110000" when sig_inp <= "00000000000001110100" else
"0100110000011001" when sig_inp <= "00000000000001110101" else
"0100101111000010" when sig_inp <= "00000000000001110110" else
"0100101101101100" when sig_inp <= "00000000000001110111" else
"0100101100010111" when sig_inp <= "00000000000001111000" else
"0100101011000001" when sig_inp <= "00000000000001111001" else
"0100101001101101" when sig_inp <= "00000000000001111010" else
"0100101000011000" when sig_inp <= "00000000000001111011" else
"0100100111000100" when sig_inp <= "00000000000001111100" else
"0100100101110000" when sig_inp <= "00000000000001111101" else
"0100100100011101" when sig_inp <= "00000000000001111110" else
"0100100011001010" when sig_inp <= "00000000000001111111" else
"0100100001110111" when sig_inp <= "00000000000010000000" else
"0100100000100101" when sig_inp <= "00000000000010000001" else
"0100011111010011" when sig_inp <= "00000000000010000010" else
"0100011110000010" when sig_inp <= "00000000000010000011" else
"0100011100110000" when sig_inp <= "00000000000010000100" else
"0100011011100000" when sig_inp <= "00000000000010000101" else
"0100011010001111" when sig_inp <= "00000000000010000110" else
"0100011000111111" when sig_inp <= "00000000000010000111" else
"0100010111101111" when sig_inp <= "00000000000010001000" else
"0100010110100000" when sig_inp <= "00000000000010001001" else
"0100010101010001" when sig_inp <= "00000000000010001010" else
"0100010100000010" when sig_inp <= "00000000000010001011" else
"0100010010110100" when sig_inp <= "00000000000010001100" else
"0100010001100110" when sig_inp <= "00000000000010001101" else
"0100010000011000" when sig_inp <= "00000000000010001110" else
"0100001111001011" when sig_inp <= "00000000000010001111" else
"0100001101111110" when sig_inp <= "00000000000010010000" else
"0100001100110001" when sig_inp <= "00000000000010010001" else
"0100001011100101" when sig_inp <= "00000000000010010010" else
"0100001010011001" when sig_inp <= "00000000000010010011" else
"0100001001001101" when sig_inp <= "00000000000010010100" else
"0100001000000010" when sig_inp <= "00000000000010010101" else
"0100000110110111" when sig_inp <= "00000000000010010110" else
"0100000101101101" when sig_inp <= "00000000000010010111" else
"0100000100100010" when sig_inp <= "00000000000010011000" else
"0100000011011000" when sig_inp <= "00000000000010011001" else
"0100000010001111" when sig_inp <= "00000000000010011010" else
"0100000001000101" when sig_inp <= "00000000000010011011" else
"0011111111111100" when sig_inp <= "00000000000010011100" else
"0011111110110100" when sig_inp <= "00000000000010011101" else
"0011111101101011" when sig_inp <= "00000000000010011110" else
"0011111100100011" when sig_inp <= "00000000000010011111" else
"0011111011011100" when sig_inp <= "00000000000010100000" else
"0011111010010100" when sig_inp <= "00000000000010100001" else
"0011111001001101" when sig_inp <= "00000000000010100010" else
"0011111000000111" when sig_inp <= "00000000000010100011" else
"0011110111000000" when sig_inp <= "00000000000010100100" else
"0011110101111010" when sig_inp <= "00000000000010100101" else
"0011110100110100" when sig_inp <= "00000000000010100110" else
"0011110011101111" when sig_inp <= "00000000000010100111" else
"0011110010101010" when sig_inp <= "00000000000010101000" else
"0011110001100101" when sig_inp <= "00000000000010101001" else
"0011110000100000" when sig_inp <= "00000000000010101010" else
"0011101111011100" when sig_inp <= "00000000000010101011" else
"0011101110011000" when sig_inp <= "00000000000010101100" else
"0011101101010100" when sig_inp <= "00000000000010101101" else
"0011101100010001" when sig_inp <= "00000000000010101110" else
"0011101011001110" when sig_inp <= "00000000000010101111" else
"0011101010001011" when sig_inp <= "00000000000010110000" else
"0011101001001001" when sig_inp <= "00000000000010110001" else
"0011101000000111" when sig_inp <= "00000000000010110010" else
"0011100111000101" when sig_inp <= "00000000000010110011" else
"0011100110000011" when sig_inp <= "00000000000010110100" else
"0011100101000010" when sig_inp <= "00000000000010110101" else
"0011100100000001" when sig_inp <= "00000000000010110110" else
"0011100011000000" when sig_inp <= "00000000000010110111" else
"0011100010000000" when sig_inp <= "00000000000010111000" else
"0011100001000000" when sig_inp <= "00000000000010111001" else
"0011100000000000" when sig_inp <= "00000000000010111010" else
"0011011111000000" when sig_inp <= "00000000000010111011" else
"0011011110000001" when sig_inp <= "00000000000010111100" else
"0011011101000010" when sig_inp <= "00000000000010111101" else
"0011011100000011" when sig_inp <= "00000000000010111110" else
"0011011011000101" when sig_inp <= "00000000000010111111" else
"0011011010000110" when sig_inp <= "00000000000011000000" else
"0011011001001001" when sig_inp <= "00000000000011000001" else
"0011011000001011" when sig_inp <= "00000000000011000010" else
"0011010111001110" when sig_inp <= "00000000000011000011" else
"0011010110010000" when sig_inp <= "00000000000011000100" else
"0011010101010100" when sig_inp <= "00000000000011000101" else
"0011010100010111" when sig_inp <= "00000000000011000110" else
"0011010011011011" when sig_inp <= "00000000000011000111" else
"0011010010011111" when sig_inp <= "00000000000011001000" else
"0011010001100011" when sig_inp <= "00000000000011001001" else
"0011010000101000" when sig_inp <= "00000000000011001010" else
"0011001111101100" when sig_inp <= "00000000000011001011" else
"0011001110110001" when sig_inp <= "00000000000011001100" else
"0011001101110111" when sig_inp <= "00000000000011001101" else
"0011001100111100" when sig_inp <= "00000000000011001110" else
"0011001100000010" when sig_inp <= "00000000000011001111" else
"0011001011001000" when sig_inp <= "00000000000011010000" else
"0011001010001111" when sig_inp <= "00000000000011010001" else
"0011001001010101" when sig_inp <= "00000000000011010010" else
"0011001000011100" when sig_inp <= "00000000000011010011" else
"0011000111100011" when sig_inp <= "00000000000011010100" else
"0011000110101011" when sig_inp <= "00000000000011010101" else
"0011000101110010" when sig_inp <= "00000000000011010110" else
"0011000100111010" when sig_inp <= "00000000000011010111" else
"0011000100000010" when sig_inp <= "00000000000011011000" else
"0011000011001010" when sig_inp <= "00000000000011011001" else
"0011000010010011" when sig_inp <= "00000000000011011010" else
"0011000001011100" when sig_inp <= "00000000000011011011" else
"0011000000100101" when sig_inp <= "00000000000011011100" else
"0010111111101110" when sig_inp <= "00000000000011011101" else
"0010111110111000" when sig_inp <= "00000000000011011110" else
"0010111110000010" when sig_inp <= "00000000000011011111" else
"0010111101001100" when sig_inp <= "00000000000011100000" else
"0010111100010110" when sig_inp <= "00000000000011100001" else
"0010111011100001" when sig_inp <= "00000000000011100010" else
"0010111010101011" when sig_inp <= "00000000000011100011" else
"0010111001110111" when sig_inp <= "00000000000011100100" else
"0010111001000010" when sig_inp <= "00000000000011100101" else
"0010111000001101" when sig_inp <= "00000000000011100110" else
"0010110111011001" when sig_inp <= "00000000000011100111" else
"0010110110100101" when sig_inp <= "00000000000011101000" else
"0010110101110001" when sig_inp <= "00000000000011101001" else
"0010110100111110" when sig_inp <= "00000000000011101010" else
"0010110100001010" when sig_inp <= "00000000000011101011" else
"0010110011010111" when sig_inp <= "00000000000011101100" else
"0010110010100100" when sig_inp <= "00000000000011101101" else
"0010110001110001" when sig_inp <= "00000000000011101110" else
"0010110000111111" when sig_inp <= "00000000000011101111" else
"0010110000001101" when sig_inp <= "00000000000011110000" else
"0010101111011011" when sig_inp <= "00000000000011110001" else
"0010101110101001" when sig_inp <= "00000000000011110010" else
"0010101101110111" when sig_inp <= "00000000000011110011" else
"0010101101000110" when sig_inp <= "00000000000011110100" else
"0010101100010101" when sig_inp <= "00000000000011110101" else
"0010101011100100" when sig_inp <= "00000000000011110110" else
"0010101010110011" when sig_inp <= "00000000000011110111" else
"0010101010000011" when sig_inp <= "00000000000011111000" else
"0010101001010011" when sig_inp <= "00000000000011111001" else
"0010101000100010" when sig_inp <= "00000000000011111010" else
"0010100111110011" when sig_inp <= "00000000000011111011" else
"0010100111000011" when sig_inp <= "00000000000011111100" else
"0010100110010100" when sig_inp <= "00000000000011111101" else
"0010100101100100" when sig_inp <= "00000000000011111110" else
"0010100100110101" when sig_inp <= "00000000000011111111" else
"0010100100000111" when sig_inp <= "00000000000100000000" else
"0010100011011000" when sig_inp <= "00000000000100000001" else
"0010100010101010" when sig_inp <= "00000000000100000010" else
"0010100001111100" when sig_inp <= "00000000000100000011" else
"0010100001001110" when sig_inp <= "00000000000100000100" else
"0010100000100000" when sig_inp <= "00000000000100000101" else
"0010011111110010" when sig_inp <= "00000000000100000110" else
"0010011111000101" when sig_inp <= "00000000000100000111" else
"0010011110011000" when sig_inp <= "00000000000100001000" else
"0010011101101011" when sig_inp <= "00000000000100001001" else
"0010011100111110" when sig_inp <= "00000000000100001010" else
"0010011100010010" when sig_inp <= "00000000000100001011" else
"0010011011100101" when sig_inp <= "00000000000100001100" else
"0010011010111001" when sig_inp <= "00000000000100001101" else
"0010011010001101" when sig_inp <= "00000000000100001110" else
"0010011001100001" when sig_inp <= "00000000000100001111" else
"0010011000110110" when sig_inp <= "00000000000100010000" else
"0010011000001010" when sig_inp <= "00000000000100010001" else
"0010010111011111" when sig_inp <= "00000000000100010010" else
"0010010110110100" when sig_inp <= "00000000000100010011" else
"0010010110001001" when sig_inp <= "00000000000100010100" else
"0010010101011111" when sig_inp <= "00000000000100010101" else
"0010010100110100" when sig_inp <= "00000000000100010110" else
"0010010100001010" when sig_inp <= "00000000000100010111" else
"0010010011100000" when sig_inp <= "00000000000100011000" else
"0010010010110110" when sig_inp <= "00000000000100011001" else
"0010010010001100" when sig_inp <= "00000000000100011010" else
"0010010001100011" when sig_inp <= "00000000000100011011" else
"0010010000111010" when sig_inp <= "00000000000100011100" else
"0010010000010001" when sig_inp <= "00000000000100011101" else
"0010001111101000" when sig_inp <= "00000000000100011110" else
"0010001110111111" when sig_inp <= "00000000000100011111" else
"0010001110010110" when sig_inp <= "00000000000100100000" else
"0010001101101110" when sig_inp <= "00000000000100100001" else
"0010001101000110" when sig_inp <= "00000000000100100010" else
"0010001100011110" when sig_inp <= "00000000000100100011" else
"0010001011110110" when sig_inp <= "00000000000100100100" else
"0010001011001110" when sig_inp <= "00000000000100100101" else
"0010001010100110" when sig_inp <= "00000000000100100110" else
"0010001001111111" when sig_inp <= "00000000000100100111" else
"0010001001011000" when sig_inp <= "00000000000100101000" else
"0010001000110001" when sig_inp <= "00000000000100101001" else
"0010001000001010" when sig_inp <= "00000000000100101010" else
"0010000111100100" when sig_inp <= "00000000000100101011" else
"0010000110111101" when sig_inp <= "00000000000100101100" else
"0010000110010111" when sig_inp <= "00000000000100101101" else
"0010000101110001" when sig_inp <= "00000000000100101110" else
"0010000101001011" when sig_inp <= "00000000000100101111" else
"0010000100100101" when sig_inp <= "00000000000100110000" else
"0010000011111111" when sig_inp <= "00000000000100110001" else
"0010000011011010" when sig_inp <= "00000000000100110010" else
"0010000010110100" when sig_inp <= "00000000000100110011" else
"0010000010001111" when sig_inp <= "00000000000100110100" else
"0010000001101010" when sig_inp <= "00000000000100110101" else
"0010000001000110" when sig_inp <= "00000000000100110110" else
"0010000000100001" when sig_inp <= "00000000000100110111" else
"0001111111111100" when sig_inp <= "00000000000100111000" else
"0001111111011000" when sig_inp <= "00000000000100111001" else
"0001111110110100" when sig_inp <= "00000000000100111010" else
"0001111110010000" when sig_inp <= "00000000000100111011" else
"0001111101101100" when sig_inp <= "00000000000100111100" else
"0001111101001000" when sig_inp <= "00000000000100111101" else
"0001111100100101" when sig_inp <= "00000000000100111110" else
"0001111100000010" when sig_inp <= "00000000000100111111" else
"0001111011011110" when sig_inp <= "00000000000101000000" else
"0001111010111011" when sig_inp <= "00000000000101000001" else
"0001111010011000" when sig_inp <= "00000000000101000010" else
"0001111001110110" when sig_inp <= "00000000000101000011" else
"0001111001010011" when sig_inp <= "00000000000101000100" else
"0001111000110001" when sig_inp <= "00000000000101000101" else
"0001111000001110" when sig_inp <= "00000000000101000110" else
"0001110111101100" when sig_inp <= "00000000000101000111" else
"0001110111001010" when sig_inp <= "00000000000101001000" else
"0001110110101001" when sig_inp <= "00000000000101001001" else
"0001110110000111" when sig_inp <= "00000000000101001010" else
"0001110101100101" when sig_inp <= "00000000000101001011" else
"0001110101000100" when sig_inp <= "00000000000101001100" else
"0001110100100011" when sig_inp <= "00000000000101001101" else
"0001110100000010" when sig_inp <= "00000000000101001110" else
"0001110011100001" when sig_inp <= "00000000000101001111" else
"0001110011000000" when sig_inp <= "00000000000101010000" else
"0001110010011111" when sig_inp <= "00000000000101010001" else
"0001110001111111" when sig_inp <= "00000000000101010010" else
"0001110001011110" when sig_inp <= "00000000000101010011" else
"0001110000111110" when sig_inp <= "00000000000101010100" else
"0001110000011110" when sig_inp <= "00000000000101010101" else
"0001101111111110" when sig_inp <= "00000000000101010110" else
"0001101111011110" when sig_inp <= "00000000000101010111" else
"0001101110111111" when sig_inp <= "00000000000101011000" else
"0001101110011111" when sig_inp <= "00000000000101011001" else
"0001101110000000" when sig_inp <= "00000000000101011010" else
"0001101101100001" when sig_inp <= "00000000000101011011" else
"0001101101000010" when sig_inp <= "00000000000101011100" else
"0001101100100011" when sig_inp <= "00000000000101011101" else
"0001101100000100" when sig_inp <= "00000000000101011110" else
"0001101011100101" when sig_inp <= "00000000000101011111" else
"0001101011000111" when sig_inp <= "00000000000101100000" else
"0001101010101000" when sig_inp <= "00000000000101100001" else
"0001101010001010" when sig_inp <= "00000000000101100010" else
"0001101001101100" when sig_inp <= "00000000000101100011" else
"0001101001001110" when sig_inp <= "00000000000101100100" else
"0001101000110000" when sig_inp <= "00000000000101100101" else
"0001101000010010" when sig_inp <= "00000000000101100110" else
"0001100111110101" when sig_inp <= "00000000000101100111" else
"0001100111010111" when sig_inp <= "00000000000101101000" else
"0001100110111010" when sig_inp <= "00000000000101101001" else
"0001100110011101" when sig_inp <= "00000000000101101010" else
"0001100110000000" when sig_inp <= "00000000000101101011" else
"0001100101100011" when sig_inp <= "00000000000101101100" else
"0001100101000110" when sig_inp <= "00000000000101101101" else
"0001100100101001" when sig_inp <= "00000000000101101110" else
"0001100100001101" when sig_inp <= "00000000000101101111" else
"0001100011110000" when sig_inp <= "00000000000101110000" else
"0001100011010100" when sig_inp <= "00000000000101110001" else
"0001100010111000" when sig_inp <= "00000000000101110010" else
"0001100010011100" when sig_inp <= "00000000000101110011" else
"0001100010000000" when sig_inp <= "00000000000101110100" else
"0001100001100100" when sig_inp <= "00000000000101110101" else
"0001100001001000" when sig_inp <= "00000000000101110110" else
"0001100000101101" when sig_inp <= "00000000000101110111" else
"0001100000010001" when sig_inp <= "00000000000101111000" else
"0001011111110110" when sig_inp <= "00000000000101111001" else
"0001011111011011" when sig_inp <= "00000000000101111010" else
"0001011111000000" when sig_inp <= "00000000000101111011" else
"0001011110100101" when sig_inp <= "00000000000101111100" else
"0001011110001010" when sig_inp <= "00000000000101111101" else
"0001011101101111" when sig_inp <= "00000000000101111110" else
"0001011101010100" when sig_inp <= "00000000000101111111" else
"0001011100111010" when sig_inp <= "00000000000110000000" else
"0001011100100000" when sig_inp <= "00000000000110000001" else
"0001011100000101" when sig_inp <= "00000000000110000010" else
"0001011011101011" when sig_inp <= "00000000000110000011" else
"0001011011010001" when sig_inp <= "00000000000110000100" else
"0001011010110111" when sig_inp <= "00000000000110000101" else
"0001011010011101" when sig_inp <= "00000000000110000110" else
"0001011010000100" when sig_inp <= "00000000000110000111" else
"0001011001101010" when sig_inp <= "00000000000110001000" else
"0001011001010001" when sig_inp <= "00000000000110001001" else
"0001011000110111" when sig_inp <= "00000000000110001010" else
"0001011000011110" when sig_inp <= "00000000000110001011" else
"0001011000000101" when sig_inp <= "00000000000110001100" else
"0001010111101100" when sig_inp <= "00000000000110001101" else
"0001010111010011" when sig_inp <= "00000000000110001110" else
"0001010110111010" when sig_inp <= "00000000000110001111" else
"0001010110100010" when sig_inp <= "00000000000110010000" else
"0001010110001001" when sig_inp <= "00000000000110010001" else
"0001010101110001" when sig_inp <= "00000000000110010010" else
"0001010101011000" when sig_inp <= "00000000000110010011" else
"0001010101000000" when sig_inp <= "00000000000110010100" else
"0001010100101000" when sig_inp <= "00000000000110010101" else
"0001010100010000" when sig_inp <= "00000000000110010110" else
"0001010011111000" when sig_inp <= "00000000000110010111" else
"0001010011100000" when sig_inp <= "00000000000110011000" else
"0001010011001001" when sig_inp <= "00000000000110011001" else
"0001010010110001" when sig_inp <= "00000000000110011010" else
"0001010010011001" when sig_inp <= "00000000000110011011" else
"0001010010000010" when sig_inp <= "00000000000110011100" else
"0001010001101011" when sig_inp <= "00000000000110011101" else
"0001010001010100" when sig_inp <= "00000000000110011110" else
"0001010000111101" when sig_inp <= "00000000000110011111" else
"0001010000100110" when sig_inp <= "00000000000110100000" else
"0001010000001111" when sig_inp <= "00000000000110100001" else
"0001001111111000" when sig_inp <= "00000000000110100010" else
"0001001111100001" when sig_inp <= "00000000000110100011" else
"0001001111001011" when sig_inp <= "00000000000110100100" else
"0001001110110100" when sig_inp <= "00000000000110100101" else
"0001001110011110" when sig_inp <= "00000000000110100110" else
"0001001110001000" when sig_inp <= "00000000000110100111" else
"0001001101110001" when sig_inp <= "00000000000110101000" else
"0001001101011011" when sig_inp <= "00000000000110101001" else
"0001001101000101" when sig_inp <= "00000000000110101010" else
"0001001100101111" when sig_inp <= "00000000000110101011" else
"0001001100011010" when sig_inp <= "00000000000110101100" else
"0001001100000100" when sig_inp <= "00000000000110101101" else
"0001001011101110" when sig_inp <= "00000000000110101110" else
"0001001011011001" when sig_inp <= "00000000000110101111" else
"0001001011000100" when sig_inp <= "00000000000110110000" else
"0001001010101110" when sig_inp <= "00000000000110110001" else
"0001001010011001" when sig_inp <= "00000000000110110010" else
"0001001010000100" when sig_inp <= "00000000000110110011" else
"0001001001101111" when sig_inp <= "00000000000110110100" else
"0001001001011010" when sig_inp <= "00000000000110110101" else
"0001001001000101" when sig_inp <= "00000000000110110110" else
"0001001000110000" when sig_inp <= "00000000000110110111" else
"0001001000011100" when sig_inp <= "00000000000110111000" else
"0001001000000111" when sig_inp <= "00000000000110111001" else
"0001000111110011" when sig_inp <= "00000000000110111010" else
"0001000111011110" when sig_inp <= "00000000000110111011" else
"0001000111001010" when sig_inp <= "00000000000110111100" else
"0001000110110110" when sig_inp <= "00000000000110111101" else
"0001000110100010" when sig_inp <= "00000000000110111110" else
"0001000110001110" when sig_inp <= "00000000000110111111" else
"0001000101111010" when sig_inp <= "00000000000111000000" else
"0001000101100110" when sig_inp <= "00000000000111000001" else
"0001000101010010" when sig_inp <= "00000000000111000010" else
"0001000100111111" when sig_inp <= "00000000000111000011" else
"0001000100101011" when sig_inp <= "00000000000111000100" else
"0001000100010111" when sig_inp <= "00000000000111000101" else
"0001000100000100" when sig_inp <= "00000000000111000110" else
"0001000011110001" when sig_inp <= "00000000000111000111" else
"0001000011011101" when sig_inp <= "00000000000111001000" else
"0001000011001010" when sig_inp <= "00000000000111001001" else
"0001000010110111" when sig_inp <= "00000000000111001010" else
"0001000010100100" when sig_inp <= "00000000000111001011" else
"0001000010010001" when sig_inp <= "00000000000111001100" else
"0001000001111111" when sig_inp <= "00000000000111001101" else
"0001000001101100" when sig_inp <= "00000000000111001110" else
"0001000001011001" when sig_inp <= "00000000000111001111" else
"0001000001000111" when sig_inp <= "00000000000111010000" else
"0001000000110100" when sig_inp <= "00000000000111010001" else
"0001000000100010" when sig_inp <= "00000000000111010010" else
"0001000000001111" when sig_inp <= "00000000000111010011" else
"0000111111111101" when sig_inp <= "00000000000111010100" else
"0000111111101011" when sig_inp <= "00000000000111010101" else
"0000111111011001" when sig_inp <= "00000000000111010110" else
"0000111111000111" when sig_inp <= "00000000000111010111" else
"0000111110110101" when sig_inp <= "00000000000111011000" else
"0000111110100011" when sig_inp <= "00000000000111011001" else
"0000111110010001" when sig_inp <= "00000000000111011010" else
"0000111110000000" when sig_inp <= "00000000000111011011" else
"0000111101101110" when sig_inp <= "00000000000111011100" else
"0000111101011101" when sig_inp <= "00000000000111011101" else
"0000111101001011" when sig_inp <= "00000000000111011110" else
"0000111100111010" when sig_inp <= "00000000000111011111" else
"0000111100101001" when sig_inp <= "00000000000111100000" else
"0000111100010111" when sig_inp <= "00000000000111100001" else
"0000111100000110" when sig_inp <= "00000000000111100010" else
"0000111011110101" when sig_inp <= "00000000000111100011" else
"0000111011100100" when sig_inp <= "00000000000111100100" else
"0000111011010011" when sig_inp <= "00000000000111100101" else
"0000111011000010" when sig_inp <= "00000000000111100110" else
"0000111010110010" when sig_inp <= "00000000000111100111" else
"0000111010100001" when sig_inp <= "00000000000111101000" else
"0000111010010000" when sig_inp <= "00000000000111101001" else
"0000111010000000" when sig_inp <= "00000000000111101010" else
"0000111001101111" when sig_inp <= "00000000000111101011" else
"0000111001011111" when sig_inp <= "00000000000111101100" else
"0000111001001111" when sig_inp <= "00000000000111101101" else
"0000111000111110" when sig_inp <= "00000000000111101110" else
"0000111000101110" when sig_inp <= "00000000000111101111" else
"0000111000011110" when sig_inp <= "00000000000111110000" else
"0000111000001110" when sig_inp <= "00000000000111110001" else
"0000110111111110" when sig_inp <= "00000000000111110010" else
"0000110111101110" when sig_inp <= "00000000000111110011" else
"0000110111011111" when sig_inp <= "00000000000111110100" else
"0000110111001111" when sig_inp <= "00000000000111110101" else
"0000110110111111" when sig_inp <= "00000000000111110110" else
"0000110110101111" when sig_inp <= "00000000000111110111" else
"0000110110100000" when sig_inp <= "00000000000111111000" else
"0000110110010000" when sig_inp <= "00000000000111111001" else
"0000110110000001" when sig_inp <= "00000000000111111010" else
"0000110101110010" when sig_inp <= "00000000000111111011" else
"0000110101100010" when sig_inp <= "00000000000111111100" else
"0000110101010011" when sig_inp <= "00000000000111111101" else
"0000110101000100" when sig_inp <= "00000000000111111110" else
"0000110100110101" when sig_inp <= "00000000000111111111" else
"0000110100100110" when sig_inp <= "00000000001000000000" else
"0000110100010111" when sig_inp <= "00000000001000000001" else
"0000110100001000" when sig_inp <= "00000000001000000010" else
"0000110011111001" when sig_inp <= "00000000001000000011" else
"0000110011101011" when sig_inp <= "00000000001000000100" else
"0000110011011100" when sig_inp <= "00000000001000000101" else
"0000110011001101" when sig_inp <= "00000000001000000110" else
"0000110010111111" when sig_inp <= "00000000001000000111" else
"0000110010110000" when sig_inp <= "00000000001000001000" else
"0000110010100010" when sig_inp <= "00000000001000001001" else
"0000110010010100" when sig_inp <= "00000000001000001010" else
"0000110010000101" when sig_inp <= "00000000001000001011" else
"0000110001110111" when sig_inp <= "00000000001000001100" else
"0000110001101001" when sig_inp <= "00000000001000001101" else
"0000110001011011" when sig_inp <= "00000000001000001110" else
"0000110001001101" when sig_inp <= "00000000001000001111" else
"0000110000111111" when sig_inp <= "00000000001000010000" else
"0000110000110001" when sig_inp <= "00000000001000010001" else
"0000110000100011" when sig_inp <= "00000000001000010010" else
"0000110000010101" when sig_inp <= "00000000001000010011" else
"0000110000001000" when sig_inp <= "00000000001000010100" else
"0000101111111010" when sig_inp <= "00000000001000010101" else
"0000101111101100" when sig_inp <= "00000000001000010110" else
"0000101111011111" when sig_inp <= "00000000001000010111" else
"0000101111010001" when sig_inp <= "00000000001000011000" else
"0000101111000100" when sig_inp <= "00000000001000011001" else
"0000101110110111" when sig_inp <= "00000000001000011010" else
"0000101110101001" when sig_inp <= "00000000001000011011" else
"0000101110011100" when sig_inp <= "00000000001000011100" else
"0000101110001111" when sig_inp <= "00000000001000011101" else
"0000101110000010" when sig_inp <= "00000000001000011110" else
"0000101101110101" when sig_inp <= "00000000001000011111" else
"0000101101101000" when sig_inp <= "00000000001000100000" else
"0000101101011011" when sig_inp <= "00000000001000100001" else
"0000101101001110" when sig_inp <= "00000000001000100010" else
"0000101101000001" when sig_inp <= "00000000001000100011" else
"0000101100110100" when sig_inp <= "00000000001000100100" else
"0000101100101000" when sig_inp <= "00000000001000100101" else
"0000101100011011" when sig_inp <= "00000000001000100110" else
"0000101100001110" when sig_inp <= "00000000001000100111" else
"0000101100000010" when sig_inp <= "00000000001000101000" else
"0000101011110101" when sig_inp <= "00000000001000101001" else
"0000101011101001" when sig_inp <= "00000000001000101010" else
"0000101011011100" when sig_inp <= "00000000001000101011" else
"0000101011010000" when sig_inp <= "00000000001000101100" else
"0000101011000100" when sig_inp <= "00000000001000101101" else
"0000101010111000" when sig_inp <= "00000000001000101110" else
"0000101010101011" when sig_inp <= "00000000001000101111" else
"0000101010011111" when sig_inp <= "00000000001000110000" else
"0000101010010011" when sig_inp <= "00000000001000110001" else
"0000101010000111" when sig_inp <= "00000000001000110010" else
"0000101001111011" when sig_inp <= "00000000001000110011" else
"0000101001101111" when sig_inp <= "00000000001000110100" else
"0000101001100100" when sig_inp <= "00000000001000110101" else
"0000101001011000" when sig_inp <= "00000000001000110110" else
"0000101001001100" when sig_inp <= "00000000001000110111" else
"0000101001000000" when sig_inp <= "00000000001000111000" else
"0000101000110101" when sig_inp <= "00000000001000111001" else
"0000101000101001" when sig_inp <= "00000000001000111010" else
"0000101000011110" when sig_inp <= "00000000001000111011" else
"0000101000010010" when sig_inp <= "00000000001000111100" else
"0000101000000111" when sig_inp <= "00000000001000111101" else
"0000100111111011" when sig_inp <= "00000000001000111110" else
"0000100111110000" when sig_inp <= "00000000001000111111" else
"0000100111100101" when sig_inp <= "00000000001001000000" else
"0000100111011001" when sig_inp <= "00000000001001000001" else
"0000100111001110" when sig_inp <= "00000000001001000010" else
"0000100111000011" when sig_inp <= "00000000001001000011" else
"0000100110111000" when sig_inp <= "00000000001001000100" else
"0000100110101101" when sig_inp <= "00000000001001000101" else
"0000100110100010" when sig_inp <= "00000000001001000110" else
"0000100110010111" when sig_inp <= "00000000001001000111" else
"0000100110001100" when sig_inp <= "00000000001001001000" else
"0000100110000001" when sig_inp <= "00000000001001001001" else
"0000100101110111" when sig_inp <= "00000000001001001010" else
"0000100101101100" when sig_inp <= "00000000001001001011" else
"0000100101100001" when sig_inp <= "00000000001001001100" else
"0000100101010110" when sig_inp <= "00000000001001001101" else
"0000100101001100" when sig_inp <= "00000000001001001110" else
"0000100101000001" when sig_inp <= "00000000001001001111" else
"0000100100110111" when sig_inp <= "00000000001001010000" else
"0000100100101100" when sig_inp <= "00000000001001010001" else
"0000100100100010" when sig_inp <= "00000000001001010010" else
"0000100100010111" when sig_inp <= "00000000001001010011" else
"0000100100001101" when sig_inp <= "00000000001001010100" else
"0000100100000011" when sig_inp <= "00000000001001010101" else
"0000100011111001" when sig_inp <= "00000000001001010110" else
"0000100011101110" when sig_inp <= "00000000001001010111" else
"0000100011100100" when sig_inp <= "00000000001001011000" else
"0000100011011010" when sig_inp <= "00000000001001011001" else
"0000100011010000" when sig_inp <= "00000000001001011010" else
"0000100011000110" when sig_inp <= "00000000001001011011" else
"0000100010111100" when sig_inp <= "00000000001001011100" else
"0000100010110010" when sig_inp <= "00000000001001011101" else
"0000100010101000" when sig_inp <= "00000000001001011110" else
"0000100010011111" when sig_inp <= "00000000001001011111" else
"0000100010010101" when sig_inp <= "00000000001001100000" else
"0000100010001011" when sig_inp <= "00000000001001100001" else
"0000100010000001" when sig_inp <= "00000000001001100010" else
"0000100001111000" when sig_inp <= "00000000001001100011" else
"0000100001101110" when sig_inp <= "00000000001001100100" else
"0000100001100101" when sig_inp <= "00000000001001100101" else
"0000100001011011" when sig_inp <= "00000000001001100110" else
"0000100001010001" when sig_inp <= "00000000001001100111" else
"0000100001001000" when sig_inp <= "00000000001001101000" else
"0000100000111111" when sig_inp <= "00000000001001101001" else
"0000100000110101" when sig_inp <= "00000000001001101010" else
"0000100000101100" when sig_inp <= "00000000001001101011" else
"0000100000100011" when sig_inp <= "00000000001001101100" else
"0000100000011001" when sig_inp <= "00000000001001101101" else
"0000100000010000" when sig_inp <= "00000000001001101110" else
"0000100000000111" when sig_inp <= "00000000001001101111" else
"0000011111111110" when sig_inp <= "00000000001001110000" else
"0000011111110101" when sig_inp <= "00000000001001110001" else
"0000011111101100" when sig_inp <= "00000000001001110010" else
"0000011111100011" when sig_inp <= "00000000001001110011" else
"0000011111011010" when sig_inp <= "00000000001001110100" else
"0000011111010001" when sig_inp <= "00000000001001110101" else
"0000011111001000" when sig_inp <= "00000000001001110110" else
"0000011110111111" when sig_inp <= "00000000001001110111" else
"0000011110110110" when sig_inp <= "00000000001001111000" else
"0000011110101110" when sig_inp <= "00000000001001111001" else
"0000011110100101" when sig_inp <= "00000000001001111010" else
"0000011110011100" when sig_inp <= "00000000001001111011" else
"0000011110010100" when sig_inp <= "00000000001001111100" else
"0000011110001011" when sig_inp <= "00000000001001111101" else
"0000011110000011" when sig_inp <= "00000000001001111110" else
"0000011101111010" when sig_inp <= "00000000001001111111" else
"0000011101110010" when sig_inp <= "00000000001010000000" else
"0000011101101001" when sig_inp <= "00000000001010000001" else
"0000011101100001" when sig_inp <= "00000000001010000010" else
"0000011101011000" when sig_inp <= "00000000001010000011" else
"0000011101010000" when sig_inp <= "00000000001010000100" else
"0000011101001000" when sig_inp <= "00000000001010000101" else
"0000011100111111" when sig_inp <= "00000000001010000110" else
"0000011100110111" when sig_inp <= "00000000001010000111" else
"0000011100101111" when sig_inp <= "00000000001010001000" else
"0000011100100111" when sig_inp <= "00000000001010001001" else
"0000011100011111" when sig_inp <= "00000000001010001010" else
"0000011100010111" when sig_inp <= "00000000001010001011" else
"0000011100001111" when sig_inp <= "00000000001010001100" else
"0000011100000110" when sig_inp <= "00000000001010001101" else
"0000011011111111" when sig_inp <= "00000000001010001110" else
"0000011011110111" when sig_inp <= "00000000001010001111" else
"0000011011101111" when sig_inp <= "00000000001010010000" else
"0000011011100111" when sig_inp <= "00000000001010010001" else
"0000011011011111" when sig_inp <= "00000000001010010010" else
"0000011011010111" when sig_inp <= "00000000001010010011" else
"0000011011001111" when sig_inp <= "00000000001010010100" else
"0000011011001000" when sig_inp <= "00000000001010010101" else
"0000011011000000" when sig_inp <= "00000000001010010110" else
"0000011010111000" when sig_inp <= "00000000001010010111" else
"0000011010110001" when sig_inp <= "00000000001010011000" else
"0000011010101001" when sig_inp <= "00000000001010011001" else
"0000011010100010" when sig_inp <= "00000000001010011010" else
"0000011010011010" when sig_inp <= "00000000001010011011" else
"0000011010010010" when sig_inp <= "00000000001010011100" else
"0000011010001011" when sig_inp <= "00000000001010011101" else
"0000011010000100" when sig_inp <= "00000000001010011110" else
"0000011001111100" when sig_inp <= "00000000001010011111" else
"0000011001110101" when sig_inp <= "00000000001010100000" else
"0000011001101101" when sig_inp <= "00000000001010100001" else
"0000011001100110" when sig_inp <= "00000000001010100010" else
"0000011001011111" when sig_inp <= "00000000001010100011" else
"0000011001011000" when sig_inp <= "00000000001010100100" else
"0000011001010000" when sig_inp <= "00000000001010100101" else
"0000011001001001" when sig_inp <= "00000000001010100110" else
"0000011001000010" when sig_inp <= "00000000001010100111" else
"0000011000111011" when sig_inp <= "00000000001010101000" else
"0000011000110100" when sig_inp <= "00000000001010101001" else
"0000011000101101" when sig_inp <= "00000000001010101010" else
"0000011000100110" when sig_inp <= "00000000001010101011" else
"0000011000011111" when sig_inp <= "00000000001010101100" else
"0000011000011000" when sig_inp <= "00000000001010101101" else
"0000011000010001" when sig_inp <= "00000000001010101110" else
"0000011000001010" when sig_inp <= "00000000001010101111" else
"0000011000000011" when sig_inp <= "00000000001010110000" else
"0000010111111101" when sig_inp <= "00000000001010110001" else
"0000010111110110" when sig_inp <= "00000000001010110010" else
"0000010111101111" when sig_inp <= "00000000001010110011" else
"0000010111101000" when sig_inp <= "00000000001010110100" else
"0000010111100001" when sig_inp <= "00000000001010110101" else
"0000010111011011" when sig_inp <= "00000000001010110110" else
"0000010111010100" when sig_inp <= "00000000001010110111" else
"0000010111001110" when sig_inp <= "00000000001010111000" else
"0000010111000111" when sig_inp <= "00000000001010111001" else
"0000010111000000" when sig_inp <= "00000000001010111010" else
"0000010110111010" when sig_inp <= "00000000001010111011" else
"0000010110110011" when sig_inp <= "00000000001010111100" else
"0000010110101101" when sig_inp <= "00000000001010111101" else
"0000010110100110" when sig_inp <= "00000000001010111110" else
"0000010110100000" when sig_inp <= "00000000001010111111" else
"0000010110011010" when sig_inp <= "00000000001011000000" else
"0000010110010011" when sig_inp <= "00000000001011000001" else
"0000010110001101" when sig_inp <= "00000000001011000010" else
"0000010110000111" when sig_inp <= "00000000001011000011" else
"0000010110000000" when sig_inp <= "00000000001011000100" else
"0000010101111010" when sig_inp <= "00000000001011000101" else
"0000010101110100" when sig_inp <= "00000000001011000110" else
"0000010101101110" when sig_inp <= "00000000001011000111" else
"0000010101101000" when sig_inp <= "00000000001011001000" else
"0000010101100001" when sig_inp <= "00000000001011001001" else
"0000010101011011" when sig_inp <= "00000000001011001010" else
"0000010101010101" when sig_inp <= "00000000001011001011" else
"0000010101001111" when sig_inp <= "00000000001011001100" else
"0000010101001001" when sig_inp <= "00000000001011001101" else
"0000010101000011" when sig_inp <= "00000000001011001110" else
"0000010100111101" when sig_inp <= "00000000001011001111" else
"0000010100110111" when sig_inp <= "00000000001011010000" else
"0000010100110001" when sig_inp <= "00000000001011010001" else
"0000010100101011" when sig_inp <= "00000000001011010010" else
"0000010100100110" when sig_inp <= "00000000001011010011" else
"0000010100100000" when sig_inp <= "00000000001011010100" else
"0000010100011010" when sig_inp <= "00000000001011010101" else
"0000010100010100" when sig_inp <= "00000000001011010110" else
"0000010100001110" when sig_inp <= "00000000001011010111" else
"0000010100001001" when sig_inp <= "00000000001011011000" else
"0000010100000011" when sig_inp <= "00000000001011011001" else
"0000010011111101" when sig_inp <= "00000000001011011010" else
"0000010011110111" when sig_inp <= "00000000001011011011" else
"0000010011110010" when sig_inp <= "00000000001011011100" else
"0000010011101100" when sig_inp <= "00000000001011011101" else
"0000010011100111" when sig_inp <= "00000000001011011110" else
"0000010011100001" when sig_inp <= "00000000001011011111" else
"0000010011011100" when sig_inp <= "00000000001011100000" else
"0000010011010110" when sig_inp <= "00000000001011100001" else
"0000010011010001" when sig_inp <= "00000000001011100010" else
"0000010011001011" when sig_inp <= "00000000001011100011" else
"0000010011000110" when sig_inp <= "00000000001011100100" else
"0000010011000000" when sig_inp <= "00000000001011100101" else
"0000010010111011" when sig_inp <= "00000000001011100110" else
"0000010010110101" when sig_inp <= "00000000001011100111" else
"0000010010110000" when sig_inp <= "00000000001011101000" else
"0000010010101011" when sig_inp <= "00000000001011101001" else
"0000010010100101" when sig_inp <= "00000000001011101010" else
"0000010010100000" when sig_inp <= "00000000001011101011" else
"0000010010011011" when sig_inp <= "00000000001011101100" else
"0000010010010110" when sig_inp <= "00000000001011101101" else
"0000010010010000" when sig_inp <= "00000000001011101110" else
"0000010010001011" when sig_inp <= "00000000001011101111" else
"0000010010000110" when sig_inp <= "00000000001011110000" else
"0000010010000001" when sig_inp <= "00000000001011110001" else
"0000010001111100" when sig_inp <= "00000000001011110010" else
"0000010001110111" when sig_inp <= "00000000001011110011" else
"0000010001110010" when sig_inp <= "00000000001011110100" else
"0000010001101101" when sig_inp <= "00000000001011110101" else
"0000010001101000" when sig_inp <= "00000000001011110110" else
"0000010001100011" when sig_inp <= "00000000001011110111" else
"0000010001011110" when sig_inp <= "00000000001011111000" else
"0000010001011001" when sig_inp <= "00000000001011111001" else
"0000010001010100" when sig_inp <= "00000000001011111010" else
"0000010001001111" when sig_inp <= "00000000001011111011" else
"0000010001001010" when sig_inp <= "00000000001011111100" else
"0000010001000101" when sig_inp <= "00000000001011111101" else
"0000010001000000" when sig_inp <= "00000000001011111110" else
"0000010000111011" when sig_inp <= "00000000001011111111" else
"0000010000110111" when sig_inp <= "00000000001100000000" else
"0000010000110010" when sig_inp <= "00000000001100000001" else
"0000010000101101" when sig_inp <= "00000000001100000010" else
"0000010000101000" when sig_inp <= "00000000001100000011" else
"0000010000100100" when sig_inp <= "00000000001100000100" else
"0000010000011111" when sig_inp <= "00000000001100000101" else
"0000010000011010" when sig_inp <= "00000000001100000110" else
"0000010000010110" when sig_inp <= "00000000001100000111" else
"0000010000010001" when sig_inp <= "00000000001100001000" else
"0000010000001100" when sig_inp <= "00000000001100001001" else
"0000010000001000" when sig_inp <= "00000000001100001010" else
"0000010000000011" when sig_inp <= "00000000001100001011" else
"0000001111111111" when sig_inp <= "00000000001100001100" else
"0000001111111010" when sig_inp <= "00000000001100001101" else
"0000001111110101" when sig_inp <= "00000000001100001110" else
"0000001111110001" when sig_inp <= "00000000001100001111" else
"0000001111101101" when sig_inp <= "00000000001100010000" else
"0000001111101000" when sig_inp <= "00000000001100010001" else
"0000001111100100" when sig_inp <= "00000000001100010010" else
"0000001111011111" when sig_inp <= "00000000001100010011" else
"0000001111011011" when sig_inp <= "00000000001100010100" else
"0000001111010110" when sig_inp <= "00000000001100010101" else
"0000001111010010" when sig_inp <= "00000000001100010110" else
"0000001111001110" when sig_inp <= "00000000001100010111" else
"0000001111001001" when sig_inp <= "00000000001100011000" else
"0000001111000101" when sig_inp <= "00000000001100011001" else
"0000001111000001" when sig_inp <= "00000000001100011010" else
"0000001110111101" when sig_inp <= "00000000001100011011" else
"0000001110111000" when sig_inp <= "00000000001100011100" else
"0000001110110100" when sig_inp <= "00000000001100011101" else
"0000001110110000" when sig_inp <= "00000000001100011110" else
"0000001110101100" when sig_inp <= "00000000001100011111" else
"0000001110101000" when sig_inp <= "00000000001100100000" else
"0000001110100011" when sig_inp <= "00000000001100100001" else
"0000001110011111" when sig_inp <= "00000000001100100010" else
"0000001110011011" when sig_inp <= "00000000001100100011" else
"0000001110010111" when sig_inp <= "00000000001100100100" else
"0000001110010011" when sig_inp <= "00000000001100100101" else
"0000001110001111" when sig_inp <= "00000000001100100110" else
"0000001110001011" when sig_inp <= "00000000001100100111" else
"0000001110000111" when sig_inp <= "00000000001100101000" else
"0000001110000011" when sig_inp <= "00000000001100101001" else
"0000001101111111" when sig_inp <= "00000000001100101010" else
"0000001101111011" when sig_inp <= "00000000001100101011" else
"0000001101110111" when sig_inp <= "00000000001100101100" else
"0000001101110011" when sig_inp <= "00000000001100101101" else
"0000001101101111" when sig_inp <= "00000000001100101110" else
"0000001101101011" when sig_inp <= "00000000001100101111" else
"0000001101100111" when sig_inp <= "00000000001100110000" else
"0000001101100011" when sig_inp <= "00000000001100110001" else
"0000001101100000" when sig_inp <= "00000000001100110010" else
"0000001101011100" when sig_inp <= "00000000001100110011" else
"0000001101011000" when sig_inp <= "00000000001100110100" else
"0000001101010100" when sig_inp <= "00000000001100110101" else
"0000001101010000" when sig_inp <= "00000000001100110110" else
"0000001101001101" when sig_inp <= "00000000001100110111" else
"0000001101001001" when sig_inp <= "00000000001100111000" else
"0000001101000101" when sig_inp <= "00000000001100111001" else
"0000001101000001" when sig_inp <= "00000000001100111010" else
"0000001100111110" when sig_inp <= "00000000001100111011" else
"0000001100111010" when sig_inp <= "00000000001100111100" else
"0000001100110110" when sig_inp <= "00000000001100111101" else
"0000001100110011" when sig_inp <= "00000000001100111110" else
"0000001100101111" when sig_inp <= "00000000001100111111" else
"0000001100101011" when sig_inp <= "00000000001101000000" else
"0000001100101000" when sig_inp <= "00000000001101000001" else
"0000001100100100" when sig_inp <= "00000000001101000010" else
"0000001100100001" when sig_inp <= "00000000001101000011" else
"0000001100011101" when sig_inp <= "00000000001101000100" else
"0000001100011010" when sig_inp <= "00000000001101000101" else
"0000001100010110" when sig_inp <= "00000000001101000110" else
"0000001100010011" when sig_inp <= "00000000001101000111" else
"0000001100001111" when sig_inp <= "00000000001101001000" else
"0000001100001100" when sig_inp <= "00000000001101001001" else
"0000001100001000" when sig_inp <= "00000000001101001010" else
"0000001100000101" when sig_inp <= "00000000001101001011" else
"0000001100000001" when sig_inp <= "00000000001101001100" else
"0000001011111110" when sig_inp <= "00000000001101001101" else
"0000001011111010" when sig_inp <= "00000000001101001110" else
"0000001011110111" when sig_inp <= "00000000001101001111" else
"0000001011110100" when sig_inp <= "00000000001101010000" else
"0000001011110000" when sig_inp <= "00000000001101010001" else
"0000001011101101" when sig_inp <= "00000000001101010010" else
"0000001011101010" when sig_inp <= "00000000001101010011" else
"0000001011100110" when sig_inp <= "00000000001101010100" else
"0000001011100011" when sig_inp <= "00000000001101010101" else
"0000001011100000" when sig_inp <= "00000000001101010110" else
"0000001011011101" when sig_inp <= "00000000001101010111" else
"0000001011011001" when sig_inp <= "00000000001101011000" else
"0000001011010110" when sig_inp <= "00000000001101011001" else
"0000001011010011" when sig_inp <= "00000000001101011010" else
"0000001011010000" when sig_inp <= "00000000001101011011" else
"0000001011001100" when sig_inp <= "00000000001101011100" else
"0000001011001001" when sig_inp <= "00000000001101011101" else
"0000001011000110" when sig_inp <= "00000000001101011110" else
"0000001011000011" when sig_inp <= "00000000001101011111" else
"0000001011000000" when sig_inp <= "00000000001101100000" else
"0000001010111101" when sig_inp <= "00000000001101100001" else
"0000001010111010" when sig_inp <= "00000000001101100010" else
"0000001010110110" when sig_inp <= "00000000001101100011" else
"0000001010110011" when sig_inp <= "00000000001101100100" else
"0000001010110000" when sig_inp <= "00000000001101100101" else
"0000001010101101" when sig_inp <= "00000000001101100110" else
"0000001010101010" when sig_inp <= "00000000001101100111" else
"0000001010100111" when sig_inp <= "00000000001101101000" else
"0000001010100100" when sig_inp <= "00000000001101101001" else
"0000001010100001" when sig_inp <= "00000000001101101010" else
"0000001010011110" when sig_inp <= "00000000001101101011" else
"0000001010011011" when sig_inp <= "00000000001101101100" else
"0000001010011000" when sig_inp <= "00000000001101101101" else
"0000001010010101" when sig_inp <= "00000000001101101110" else
"0000001010010010" when sig_inp <= "00000000001101101111" else
"0000001010001111" when sig_inp <= "00000000001101110000" else
"0000001010001101" when sig_inp <= "00000000001101110001" else
"0000001010001010" when sig_inp <= "00000000001101110010" else
"0000001010000111" when sig_inp <= "00000000001101110011" else
"0000001010000100" when sig_inp <= "00000000001101110100" else
"0000001010000001" when sig_inp <= "00000000001101110101" else
"0000001001111110" when sig_inp <= "00000000001101110110" else
"0000001001111011" when sig_inp <= "00000000001101110111" else
"0000001001111001" when sig_inp <= "00000000001101111000" else
"0000001001110110" when sig_inp <= "00000000001101111001" else
"0000001001110011" when sig_inp <= "00000000001101111010" else
"0000001001110000" when sig_inp <= "00000000001101111011" else
"0000001001101101" when sig_inp <= "00000000001101111100" else
"0000001001101011" when sig_inp <= "00000000001101111101" else
"0000001001101000" when sig_inp <= "00000000001101111110" else
"0000001001100101" when sig_inp <= "00000000001101111111" else
"0000001001100010" when sig_inp <= "00000000001110000000" else
"0000001001100000" when sig_inp <= "00000000001110000001" else
"0000001001011101" when sig_inp <= "00000000001110000010" else
"0000001001011010" when sig_inp <= "00000000001110000011" else
"0000001001011000" when sig_inp <= "00000000001110000100" else
"0000001001010101" when sig_inp <= "00000000001110000101" else
"0000001001010010" when sig_inp <= "00000000001110000110" else
"0000001001010000" when sig_inp <= "00000000001110000111" else
"0000001001001101" when sig_inp <= "00000000001110001000" else
"0000001001001010" when sig_inp <= "00000000001110001001" else
"0000001001001000" when sig_inp <= "00000000001110001010" else
"0000001001000101" when sig_inp <= "00000000001110001011" else
"0000001001000011" when sig_inp <= "00000000001110001100" else
"0000001001000000" when sig_inp <= "00000000001110001101" else
"0000001000111110" when sig_inp <= "00000000001110001110" else
"0000001000111011" when sig_inp <= "00000000001110001111" else
"0000001000111000" when sig_inp <= "00000000001110010000" else
"0000001000110110" when sig_inp <= "00000000001110010001" else
"0000001000110011" when sig_inp <= "00000000001110010010" else
"0000001000110001" when sig_inp <= "00000000001110010011" else
"0000001000101110" when sig_inp <= "00000000001110010100" else
"0000001000101100" when sig_inp <= "00000000001110010101" else
"0000001000101010" when sig_inp <= "00000000001110010110" else
"0000001000100111" when sig_inp <= "00000000001110010111" else
"0000001000100101" when sig_inp <= "00000000001110011000" else
"0000001000100010" when sig_inp <= "00000000001110011001" else
"0000001000100000" when sig_inp <= "00000000001110011010" else
"0000001000011101" when sig_inp <= "00000000001110011011" else
"0000001000011011" when sig_inp <= "00000000001110011100" else
"0000001000011001" when sig_inp <= "00000000001110011101" else
"0000001000010110" when sig_inp <= "00000000001110011110" else
"0000001000010100" when sig_inp <= "00000000001110011111" else
"0000001000010001" when sig_inp <= "00000000001110100000" else
"0000001000001111" when sig_inp <= "00000000001110100001" else
"0000001000001101" when sig_inp <= "00000000001110100010" else
"0000001000001010" when sig_inp <= "00000000001110100011" else
"0000001000001000" when sig_inp <= "00000000001110100100" else
"0000001000000110" when sig_inp <= "00000000001110100101" else
"0000001000000011" when sig_inp <= "00000000001110100110" else
"0000001000000001" when sig_inp <= "00000000001110100111" else
"0000000111111111" when sig_inp <= "00000000001110101000" else
"0000000111111101" when sig_inp <= "00000000001110101001" else
"0000000111111010" when sig_inp <= "00000000001110101010" else
"0000000111111000" when sig_inp <= "00000000001110101011" else
"0000000111110110" when sig_inp <= "00000000001110101100" else
"0000000111110100" when sig_inp <= "00000000001110101101" else
"0000000111110001" when sig_inp <= "00000000001110101110" else
"0000000111101111" when sig_inp <= "00000000001110101111" else
"0000000111101101" when sig_inp <= "00000000001110110000" else
"0000000111101011" when sig_inp <= "00000000001110110001" else
"0000000111101001" when sig_inp <= "00000000001110110010" else
"0000000111100111" when sig_inp <= "00000000001110110011" else
"0000000111100100" when sig_inp <= "00000000001110110100" else
"0000000111100010" when sig_inp <= "00000000001110110101" else
"0000000111100000" when sig_inp <= "00000000001110110110" else
"0000000111011110" when sig_inp <= "00000000001110110111" else
"0000000111011100" when sig_inp <= "00000000001110111000" else
"0000000111011010" when sig_inp <= "00000000001110111001" else
"0000000111011000" when sig_inp <= "00000000001110111010" else
"0000000111010110" when sig_inp <= "00000000001110111011" else
"0000000111010011" when sig_inp <= "00000000001110111100" else
"0000000111010001" when sig_inp <= "00000000001110111101" else
"0000000111001111" when sig_inp <= "00000000001110111110" else
"0000000111001101" when sig_inp <= "00000000001110111111" else
"0000000111001011" when sig_inp <= "00000000001111000000" else
"0000000111001001" when sig_inp <= "00000000001111000001" else
"0000000111000111" when sig_inp <= "00000000001111000010" else
"0000000111000101" when sig_inp <= "00000000001111000011" else
"0000000111000011" when sig_inp <= "00000000001111000100" else
"0000000111000001" when sig_inp <= "00000000001111000101" else
"0000000110111111" when sig_inp <= "00000000001111000110" else
"0000000110111101" when sig_inp <= "00000000001111000111" else
"0000000110111011" when sig_inp <= "00000000001111001000" else
"0000000110111001" when sig_inp <= "00000000001111001001" else
"0000000110110111" when sig_inp <= "00000000001111001010" else
"0000000110110101" when sig_inp <= "00000000001111001011" else
"0000000110110011" when sig_inp <= "00000000001111001100" else
"0000000110110001" when sig_inp <= "00000000001111001101" else
"0000000110101111" when sig_inp <= "00000000001111001110" else
"0000000110101110" when sig_inp <= "00000000001111001111" else
"0000000110101100" when sig_inp <= "00000000001111010000" else
"0000000110101010" when sig_inp <= "00000000001111010001" else
"0000000110101000" when sig_inp <= "00000000001111010010" else
"0000000110100110" when sig_inp <= "00000000001111010011" else
"0000000110100100" when sig_inp <= "00000000001111010100" else
"0000000110100010" when sig_inp <= "00000000001111010101" else
"0000000110100000" when sig_inp <= "00000000001111010110" else
"0000000110011111" when sig_inp <= "00000000001111010111" else
"0000000110011101" when sig_inp <= "00000000001111011000" else
"0000000110011011" when sig_inp <= "00000000001111011001" else
"0000000110011001" when sig_inp <= "00000000001111011010" else
"0000000110010111" when sig_inp <= "00000000001111011011" else
"0000000110010101" when sig_inp <= "00000000001111011100" else
"0000000110010100" when sig_inp <= "00000000001111011101" else
"0000000110010010" when sig_inp <= "00000000001111011110" else
"0000000110010000" when sig_inp <= "00000000001111011111" else
"0000000110001110" when sig_inp <= "00000000001111100000" else
"0000000110001100" when sig_inp <= "00000000001111100001" else
"0000000110001011" when sig_inp <= "00000000001111100010" else
"0000000110001001" when sig_inp <= "00000000001111100011" else
"0000000110000111" when sig_inp <= "00000000001111100100" else
"0000000110000101" when sig_inp <= "00000000001111100101" else
"0000000110000100" when sig_inp <= "00000000001111100110" else
"0000000110000010" when sig_inp <= "00000000001111100111" else
"0000000110000000" when sig_inp <= "00000000001111101000" else
"0000000101111111" when sig_inp <= "00000000001111101001" else
"0000000101111101" when sig_inp <= "00000000001111101010" else
"0000000101111011" when sig_inp <= "00000000001111101011" else
"0000000101111010" when sig_inp <= "00000000001111101100" else
"0000000101111000" when sig_inp <= "00000000001111101101" else
"0000000101110110" when sig_inp <= "00000000001111101110" else
"0000000101110101" when sig_inp <= "00000000001111101111" else
"0000000101110011" when sig_inp <= "00000000001111110000" else
"0000000101110001" when sig_inp <= "00000000001111110001" else
"0000000101110000" when sig_inp <= "00000000001111110010" else
"0000000101101110" when sig_inp <= "00000000001111110011" else
"0000000101101100" when sig_inp <= "00000000001111110100" else
"0000000101101011" when sig_inp <= "00000000001111110101" else
"0000000101101001" when sig_inp <= "00000000001111110110" else
"0000000101100111" when sig_inp <= "00000000001111110111" else
"0000000101100110" when sig_inp <= "00000000001111111000" else
"0000000101100100" when sig_inp <= "00000000001111111001" else
"0000000101100011" when sig_inp <= "00000000001111111010" else
"0000000101100001" when sig_inp <= "00000000001111111011" else
"0000000101100000" when sig_inp <= "00000000001111111100" else
"0000000101011110" when sig_inp <= "00000000001111111101" else
"0000000101011100" when sig_inp <= "00000000001111111110" else
"0000000101011011" when sig_inp <= "00000000001111111111" else
"0000000101011001" when sig_inp <= "00000000010000000000" else
"0000000101011000" when sig_inp <= "00000000010000000001" else
"0000000101010110" when sig_inp <= "00000000010000000010" else
"0000000101010101" when sig_inp <= "00000000010000000011" else
"0000000101010011" when sig_inp <= "00000000010000000100" else
"0000000101010010" when sig_inp <= "00000000010000000101" else
"0000000101010000" when sig_inp <= "00000000010000000110" else
"0000000101001111" when sig_inp <= "00000000010000000111" else
"0000000101001101" when sig_inp <= "00000000010000001000" else
"0000000101001100" when sig_inp <= "00000000010000001001" else
"0000000101001010" when sig_inp <= "00000000010000001010" else
"0000000101001001" when sig_inp <= "00000000010000001011" else
"0000000101000111" when sig_inp <= "00000000010000001100" else
"0000000101000110" when sig_inp <= "00000000010000001101" else
"0000000101000101" when sig_inp <= "00000000010000001110" else
"0000000101000011" when sig_inp <= "00000000010000001111" else
"0000000101000010" when sig_inp <= "00000000010000010000" else
"0000000101000000" when sig_inp <= "00000000010000010001" else
"0000000100111111" when sig_inp <= "00000000010000010010" else
"0000000100111101" when sig_inp <= "00000000010000010011" else
"0000000100111100" when sig_inp <= "00000000010000010100" else
"0000000100111011" when sig_inp <= "00000000010000010101" else
"0000000100111001" when sig_inp <= "00000000010000010110" else
"0000000100111000" when sig_inp <= "00000000010000010111" else
"0000000100110110" when sig_inp <= "00000000010000011000" else
"0000000100110101" when sig_inp <= "00000000010000011001" else
"0000000100110100" when sig_inp <= "00000000010000011010" else
"0000000100110010" when sig_inp <= "00000000010000011011" else
"0000000100110001" when sig_inp <= "00000000010000011100" else
"0000000100110000" when sig_inp <= "00000000010000011101" else
"0000000100101110" when sig_inp <= "00000000010000011110" else
"0000000100101101" when sig_inp <= "00000000010000011111" else
"0000000100101100" when sig_inp <= "00000000010000100000" else
"0000000100101010" when sig_inp <= "00000000010000100001" else
"0000000100101001" when sig_inp <= "00000000010000100010" else
"0000000100101000" when sig_inp <= "00000000010000100011" else
"0000000100100110" when sig_inp <= "00000000010000100100" else
"0000000100100101" when sig_inp <= "00000000010000100101" else
"0000000100100100" when sig_inp <= "00000000010000100110" else
"0000000100100010" when sig_inp <= "00000000010000100111" else
"0000000100100001" when sig_inp <= "00000000010000101000" else
"0000000100100000" when sig_inp <= "00000000010000101001" else
"0000000100011110" when sig_inp <= "00000000010000101010" else
"0000000100011101" when sig_inp <= "00000000010000101011" else
"0000000100011100" when sig_inp <= "00000000010000101100" else
"0000000100011011" when sig_inp <= "00000000010000101101" else
"0000000100011001" when sig_inp <= "00000000010000101110" else
"0000000100011000" when sig_inp <= "00000000010000101111" else
"0000000100010111" when sig_inp <= "00000000010000110000" else
"0000000100010110" when sig_inp <= "00000000010000110001" else
"0000000100010100" when sig_inp <= "00000000010000110010" else
"0000000100010011" when sig_inp <= "00000000010000110011" else
"0000000100010010" when sig_inp <= "00000000010000110100" else
"0000000100010001" when sig_inp <= "00000000010000110101" else
"0000000100010000" when sig_inp <= "00000000010000110110" else
"0000000100001110" when sig_inp <= "00000000010000110111" else
"0000000100001101" when sig_inp <= "00000000010000111000" else
"0000000100001100" when sig_inp <= "00000000010000111001" else
"0000000100001011" when sig_inp <= "00000000010000111010" else
"0000000100001010" when sig_inp <= "00000000010000111011" else
"0000000100001000" when sig_inp <= "00000000010000111100" else
"0000000100000111" when sig_inp <= "00000000010000111101" else
"0000000100000110" when sig_inp <= "00000000010000111110" else
"0000000100000101" when sig_inp <= "00000000010000111111" else
"0000000100000100" when sig_inp <= "00000000010001000000" else
"0000000100000011" when sig_inp <= "00000000010001000001" else
"0000000100000001" when sig_inp <= "00000000010001000010" else
"0000000100000000" when sig_inp <= "00000000010001000011" else
"0000000011111111" when sig_inp <= "00000000010001000100" else
"0000000011111110" when sig_inp <= "00000000010001000101" else
"0000000011111101" when sig_inp <= "00000000010001000110" else
"0000000011111100" when sig_inp <= "00000000010001000111" else
"0000000011111011" when sig_inp <= "00000000010001001000" else
"0000000011111010" when sig_inp <= "00000000010001001001" else
"0000000011111000" when sig_inp <= "00000000010001001010" else
"0000000011110111" when sig_inp <= "00000000010001001011" else
"0000000011110110" when sig_inp <= "00000000010001001100" else
"0000000011110101" when sig_inp <= "00000000010001001101" else
"0000000011110100" when sig_inp <= "00000000010001001110" else
"0000000011110011" when sig_inp <= "00000000010001001111" else
"0000000011110010" when sig_inp <= "00000000010001010000" else
"0000000011110001" when sig_inp <= "00000000010001010001" else
"0000000011110000" when sig_inp <= "00000000010001010010" else
"0000000011101111" when sig_inp <= "00000000010001010011" else
"0000000011101110" when sig_inp <= "00000000010001010100" else
"0000000011101101" when sig_inp <= "00000000010001010101" else
"0000000011101100" when sig_inp <= "00000000010001010110" else
"0000000011101010" when sig_inp <= "00000000010001010111" else
"0000000011101001" when sig_inp <= "00000000010001011000" else
"0000000011101000" when sig_inp <= "00000000010001011001" else
"0000000011100111" when sig_inp <= "00000000010001011010" else
"0000000011100110" when sig_inp <= "00000000010001011011" else
"0000000011100101" when sig_inp <= "00000000010001011100" else
"0000000011100100" when sig_inp <= "00000000010001011101" else
"0000000011100011" when sig_inp <= "00000000010001011110" else
"0000000011100010" when sig_inp <= "00000000010001011111" else
"0000000011100001" when sig_inp <= "00000000010001100000" else
"0000000011100000" when sig_inp <= "00000000010001100001" else
"0000000011011111" when sig_inp <= "00000000010001100010" else
"0000000011011110" when sig_inp <= "00000000010001100011" else
"0000000011011101" when sig_inp <= "00000000010001100100" else
"0000000011011100" when sig_inp <= "00000000010001100101" else
"0000000011011011" when sig_inp <= "00000000010001100110" else
"0000000011011010" when sig_inp <= "00000000010001100111" else
"0000000011011001" when sig_inp <= "00000000010001101000" else
"0000000011011000" when sig_inp <= "00000000010001101001" else
"0000000011010111" when sig_inp <= "00000000010001101010" else
"0000000011010110" when sig_inp <= "00000000010001101011" else
"0000000011010101" when sig_inp <= "00000000010001101101" else
"0000000011010100" when sig_inp <= "00000000010001101110" else
"0000000011010011" when sig_inp <= "00000000010001101111" else
"0000000011010010" when sig_inp <= "00000000010001110000" else
"0000000011010001" when sig_inp <= "00000000010001110001" else
"0000000011010000" when sig_inp <= "00000000010001110010" else
"0000000011001111" when sig_inp <= "00000000010001110011" else
"0000000011001110" when sig_inp <= "00000000010001110100" else
"0000000011001101" when sig_inp <= "00000000010001110101" else
"0000000011001100" when sig_inp <= "00000000010001110110" else
"0000000011001011" when sig_inp <= "00000000010001110111" else
"0000000011001010" when sig_inp <= "00000000010001111000" else
"0000000011001001" when sig_inp <= "00000000010001111010" else
"0000000011001000" when sig_inp <= "00000000010001111011" else
"0000000011000111" when sig_inp <= "00000000010001111100" else
"0000000011000110" when sig_inp <= "00000000010001111101" else
"0000000011000101" when sig_inp <= "00000000010001111110" else
"0000000011000100" when sig_inp <= "00000000010001111111" else
"0000000011000011" when sig_inp <= "00000000010010000000" else
"0000000011000010" when sig_inp <= "00000000010010000001" else
"0000000011000001" when sig_inp <= "00000000010010000011" else
"0000000011000000" when sig_inp <= "00000000010010000100" else
"0000000010111111" when sig_inp <= "00000000010010000101" else
"0000000010111110" when sig_inp <= "00000000010010000110" else
"0000000010111101" when sig_inp <= "00000000010010000111" else
"0000000010111100" when sig_inp <= "00000000010010001000" else
"0000000010111011" when sig_inp <= "00000000010010001010" else
"0000000010111010" when sig_inp <= "00000000010010001011" else
"0000000010111001" when sig_inp <= "00000000010010001100" else
"0000000010111000" when sig_inp <= "00000000010010001101" else
"0000000010110111" when sig_inp <= "00000000010010001111" else
"0000000010110110" when sig_inp <= "00000000010010010000" else
"0000000010110101" when sig_inp <= "00000000010010010001" else
"0000000010110100" when sig_inp <= "00000000010010010010" else
"0000000010110011" when sig_inp <= "00000000010010010011" else
"0000000010110010" when sig_inp <= "00000000010010010101" else
"0000000010110001" when sig_inp <= "00000000010010010110" else
"0000000010110000" when sig_inp <= "00000000010010010111" else
"0000000010101111" when sig_inp <= "00000000010010011001" else
"0000000010101110" when sig_inp <= "00000000010010011010" else
"0000000010101101" when sig_inp <= "00000000010010011011" else
"0000000010101100" when sig_inp <= "00000000010010011100" else
"0000000010101011" when sig_inp <= "00000000010010011110" else
"0000000010101010" when sig_inp <= "00000000010010011111" else
"0000000010101001" when sig_inp <= "00000000010010100000" else
"0000000010101000" when sig_inp <= "00000000010010100010" else
"0000000010100111" when sig_inp <= "00000000010010100011" else
"0000000010100110" when sig_inp <= "00000000010010100100" else
"0000000010100101" when sig_inp <= "00000000010010100110" else
"0000000010100100" when sig_inp <= "00000000010010100111" else
"0000000010100011" when sig_inp <= "00000000010010101000" else
"0000000010100010" when sig_inp <= "00000000010010101010" else
"0000000010100001" when sig_inp <= "00000000010010101011" else
"0000000010100000" when sig_inp <= "00000000010010101101" else
"0000000010011111" when sig_inp <= "00000000010010101110" else
"0000000010011110" when sig_inp <= "00000000010010101111" else
"0000000010011101" when sig_inp <= "00000000010010110001" else
"0000000010011100" when sig_inp <= "00000000010010110010" else
"0000000010011011" when sig_inp <= "00000000010010110100" else
"0000000010011010" when sig_inp <= "00000000010010110101" else
"0000000010011001" when sig_inp <= "00000000010010110111" else
"0000000010011000" when sig_inp <= "00000000010010111000" else
"0000000010010111" when sig_inp <= "00000000010010111001" else
"0000000010010110" when sig_inp <= "00000000010010111011" else
"0000000010010101" when sig_inp <= "00000000010010111100" else
"0000000010010100" when sig_inp <= "00000000010010111110" else
"0000000010010011" when sig_inp <= "00000000010010111111" else
"0000000010010010" when sig_inp <= "00000000010011000001" else
"0000000010010001" when sig_inp <= "00000000010011000011" else
"0000000010010000" when sig_inp <= "00000000010011000100" else
"0000000010001111" when sig_inp <= "00000000010011000110" else
"0000000010001110" when sig_inp <= "00000000010011000111" else
"0000000010001101" when sig_inp <= "00000000010011001001" else
"0000000010001100" when sig_inp <= "00000000010011001010" else
"0000000010001011" when sig_inp <= "00000000010011001100" else
"0000000010001010" when sig_inp <= "00000000010011001110" else
"0000000010001001" when sig_inp <= "00000000010011001111" else
"0000000010001000" when sig_inp <= "00000000010011010001" else
"0000000010000111" when sig_inp <= "00000000010011010011" else
"0000000010000110" when sig_inp <= "00000000010011010100" else
"0000000010000101" when sig_inp <= "00000000010011010110" else
"0000000010000100" when sig_inp <= "00000000010011011000" else
"0000000010000011" when sig_inp <= "00000000010011011001" else
"0000000010000010" when sig_inp <= "00000000010011011011" else
"0000000010000001" when sig_inp <= "00000000010011011101" else
"0000000010000000" when sig_inp <= "00000000010011011110" else
"0000000001111111" when sig_inp <= "00000000010011100000" else
"0000000001111110" when sig_inp <= "00000000010011100010" else
"0000000001111101" when sig_inp <= "00000000010011100100" else
"0000000001111100" when sig_inp <= "00000000010011100110" else
"0000000001111011" when sig_inp <= "00000000010011100111" else
"0000000001111010" when sig_inp <= "00000000010011101001" else
"0000000001111001" when sig_inp <= "00000000010011101011" else
"0000000001111000" when sig_inp <= "00000000010011101101" else
"0000000001110111" when sig_inp <= "00000000010011101111" else
"0000000001110110" when sig_inp <= "00000000010011110001" else
"0000000001110101" when sig_inp <= "00000000010011110010" else
"0000000001110100" when sig_inp <= "00000000010011110100" else
"0000000001110011" when sig_inp <= "00000000010011110110" else
"0000000001110010" when sig_inp <= "00000000010011111000" else
"0000000001110001" when sig_inp <= "00000000010011111010" else
"0000000001110000" when sig_inp <= "00000000010011111100" else
"0000000001101111" when sig_inp <= "00000000010011111110" else
"0000000001101110" when sig_inp <= "00000000010100000000" else
"0000000001101101" when sig_inp <= "00000000010100000010" else
"0000000001101100" when sig_inp <= "00000000010100000100" else
"0000000001101011" when sig_inp <= "00000000010100000110" else
"0000000001101010" when sig_inp <= "00000000010100001000" else
"0000000001101001" when sig_inp <= "00000000010100001011" else
"0000000001101000" when sig_inp <= "00000000010100001101" else
"0000000001100111" when sig_inp <= "00000000010100001111" else
"0000000001100110" when sig_inp <= "00000000010100010001" else
"0000000001100101" when sig_inp <= "00000000010100010011" else
"0000000001100100" when sig_inp <= "00000000010100010101" else
"0000000001100011" when sig_inp <= "00000000010100011000" else
"0000000001100010" when sig_inp <= "00000000010100011010" else
"0000000001100001" when sig_inp <= "00000000010100011100" else
"0000000001100000" when sig_inp <= "00000000010100011111" else
"0000000001011111" when sig_inp <= "00000000010100100001" else
"0000000001011110" when sig_inp <= "00000000010100100011" else
"0000000001011101" when sig_inp <= "00000000010100100110" else
"0000000001011100" when sig_inp <= "00000000010100101000" else
"0000000001011011" when sig_inp <= "00000000010100101010" else
"0000000001011010" when sig_inp <= "00000000010100101101" else
"0000000001011001" when sig_inp <= "00000000010100101111" else
"0000000001011000" when sig_inp <= "00000000010100110010" else
"0000000001010111" when sig_inp <= "00000000010100110100" else
"0000000001010110" when sig_inp <= "00000000010100110111" else
"0000000001010101" when sig_inp <= "00000000010100111010" else
"0000000001010100" when sig_inp <= "00000000010100111100" else
"0000000001010011" when sig_inp <= "00000000010100111111" else
"0000000001010010" when sig_inp <= "00000000010101000010" else
"0000000001010001" when sig_inp <= "00000000010101000100" else
"0000000001010000" when sig_inp <= "00000000010101000111" else
"0000000001001111" when sig_inp <= "00000000010101001010" else
"0000000001001110" when sig_inp <= "00000000010101001101" else
"0000000001001101" when sig_inp <= "00000000010101010000" else
"0000000001001100" when sig_inp <= "00000000010101010011" else
"0000000001001011" when sig_inp <= "00000000010101010101" else
"0000000001001010" when sig_inp <= "00000000010101011000" else
"0000000001001001" when sig_inp <= "00000000010101011011" else
"0000000001001000" when sig_inp <= "00000000010101011111" else
"0000000001000111" when sig_inp <= "00000000010101100010" else
"0000000001000110" when sig_inp <= "00000000010101100101" else
"0000000001000101" when sig_inp <= "00000000010101101000" else
"0000000001000100" when sig_inp <= "00000000010101101011" else
"0000000001000011" when sig_inp <= "00000000010101101110" else
"0000000001000010" when sig_inp <= "00000000010101110010" else
"0000000001000001" when sig_inp <= "00000000010101110101" else
"0000000001000000" when sig_inp <= "00000000010101111001" else
"0000000000111111" when sig_inp <= "00000000010101111100" else
"0000000000111110" when sig_inp <= "00000000010110000000" else
"0000000000111101" when sig_inp <= "00000000010110000011" else
"0000000000111100" when sig_inp <= "00000000010110000111" else
"0000000000111011" when sig_inp <= "00000000010110001011" else
"0000000000111010" when sig_inp <= "00000000010110001110" else
"0000000000111001" when sig_inp <= "00000000010110010010" else
"0000000000111000" when sig_inp <= "00000000010110010110" else
"0000000000110111" when sig_inp <= "00000000010110011010" else
"0000000000110110" when sig_inp <= "00000000010110011110" else
"0000000000110101" when sig_inp <= "00000000010110100010" else
"0000000000110100" when sig_inp <= "00000000010110100111" else
"0000000000110011" when sig_inp <= "00000000010110101011" else
"0000000000110010" when sig_inp <= "00000000010110101111" else
"0000000000110001" when sig_inp <= "00000000010110110100" else
"0000000000110000" when sig_inp <= "00000000010110111000" else
"0000000000101111" when sig_inp <= "00000000010110111101" else
"0000000000101110" when sig_inp <= "00000000010111000010" else
"0000000000101101" when sig_inp <= "00000000010111000110" else
"0000000000101100" when sig_inp <= "00000000010111001011" else
"0000000000101011" when sig_inp <= "00000000010111010000" else
"0000000000101010" when sig_inp <= "00000000010111010110" else
"0000000000101001" when sig_inp <= "00000000010111011011" else
"0000000000101000" when sig_inp <= "00000000010111100000" else
"0000000000100111" when sig_inp <= "00000000010111100110" else
"0000000000100110" when sig_inp <= "00000000010111101100" else
"0000000000100101" when sig_inp <= "00000000010111110001" else
"0000000000100100" when sig_inp <= "00000000010111110111" else
"0000000000100011" when sig_inp <= "00000000010111111110" else
"0000000000100010" when sig_inp <= "00000000011000000100" else
"0000000000100001" when sig_inp <= "00000000011000001010" else
"0000000000100000" when sig_inp <= "00000000011000010001" else
"0000000000011111" when sig_inp <= "00000000011000011000" else
"0000000000011110" when sig_inp <= "00000000011000011111" else
"0000000000011101" when sig_inp <= "00000000011000100111" else
"0000000000011100" when sig_inp <= "00000000011000101110" else
"0000000000011011" when sig_inp <= "00000000011000110110" else
"0000000000011010" when sig_inp <= "00000000011000111110" else
"0000000000011001" when sig_inp <= "00000000011001000111" else
"0000000000011000" when sig_inp <= "00000000011001010000" else
"0000000000010111" when sig_inp <= "00000000011001011001" else
"0000000000010110" when sig_inp <= "00000000011001100010" else
"0000000000010101" when sig_inp <= "00000000011001101100" else
"0000000000010100" when sig_inp <= "00000000011001110111" else
"0000000000010011" when sig_inp <= "00000000011010000010" else
"0000000000010010" when sig_inp <= "00000000011010001101" else
"0000000000010001" when sig_inp <= "00000000011010011010" else
"0000000000010000" when sig_inp <= "00000000011010100110" else
"0000000000001111" when sig_inp <= "00000000011010110100" else
"0000000000001110" when sig_inp <= "00000000011011000011" else
"0000000000001101" when sig_inp <= "00000000011011010010" else
"0000000000001100" when sig_inp <= "00000000011011100011" else
"0000000000001011" when sig_inp <= "00000000011011110101" else
"0000000000001010" when sig_inp <= "00000000011100001000" else
"0000000000001001" when sig_inp <= "00000000011100011110" else
"0000000000001000" when sig_inp <= "00000000011100110101" else
"0000000000000111" when sig_inp <= "00000000011101010000" else
"0000000000000110" when sig_inp <= "00000000011101101110" else
"0000000000000101" when sig_inp <= "00000000011110010001" else
"0000000000000100" when sig_inp <= "00000000011110111010" else
"0000000000000011" when sig_inp <= "00000000011111101100" else
"0000000000000010" when sig_inp <= "00000000100000101101" else
"0000000000000001" when sig_inp <= "00000000100010001000" else
"0000000000000000" when sig_inp <= "00000000100100100100" else
"0000000000000000";



----------------
--"Sigma_r = 5"
--"a = 3"
-----------------------------
--"1000000000000000" when sig_inp <= "000000000000000000000000000000000000" else
--"0111111101101110" when sig_inp <= "000000000000000000000000000010010001" else
--"0111111011011110" when sig_inp <= "000000000000000000000000000100100011" else
--"0111111001001101" when sig_inp <= "000000000000000000000000000110110100" else
--"0111110110111110" when sig_inp <= "000000000000000000000000001001000110" else
--"0111110100101111" when sig_inp <= "000000000000000000000000001011011000" else
--"0111110010100001" when sig_inp <= "000000000000000000000000001101101001" else
--"0111110000010100" when sig_inp <= "000000000000000000000000001111111011" else
--"0111101110000111" when sig_inp <= "000000000000000000000000010010001101" else
--"0111101011111011" when sig_inp <= "000000000000000000000000010100011110" else
--"0111101001101111" when sig_inp <= "000000000000000000000000010110110000" else
--"0111100111100100" when sig_inp <= "000000000000000000000000011001000001" else
--"0111100101011010" when sig_inp <= "000000000000000000000000011011010011" else
--"0111100011010000" when sig_inp <= "000000000000000000000000011101100101" else
--"0111100001000111" when sig_inp <= "000000000000000000000000011111110110" else
--"0111011110111110" when sig_inp <= "000000000000000000000000100010001000" else
--"0111011100110110" when sig_inp <= "000000000000000000000000100100011010" else
--"0111011010101111" when sig_inp <= "000000000000000000000000100110101011" else
--"0111011000101000" when sig_inp <= "000000000000000000000000101000111101" else
--"0111010110100010" when sig_inp <= "000000000000000000000000101011001111" else
--"0111010100011100" when sig_inp <= "000000000000000000000000101101100000" else
--"0111010010011000" when sig_inp <= "000000000000000000000000101111110010" else
--"0111010000010011" when sig_inp <= "000000000000000000000000110010000011" else
--"0111001110001111" when sig_inp <= "000000000000000000000000110100010101" else
--"0111001100001100" when sig_inp <= "000000000000000000000000110110100111" else
--"0111001010001010" when sig_inp <= "000000000000000000000000111000111000" else
--"0111001000001000" when sig_inp <= "000000000000000000000000111011001010" else
--"0111000110000110" when sig_inp <= "000000000000000000000000111101011100" else
--"0111000100000101" when sig_inp <= "000000000000000000000000111111101101" else
--"0111000010000101" when sig_inp <= "000000000000000000000001000001111111" else
--"0111000000000101" when sig_inp <= "000000000000000000000001000100010001" else
--"0110111110000110" when sig_inp <= "000000000000000000000001000110100010" else
--"0110111100000111" when sig_inp <= "000000000000000000000001001000110100" else
--"0110111010001001" when sig_inp <= "000000000000000000000001001011000101" else
--"0110111000001100" when sig_inp <= "000000000000000000000001001101010111" else
--"0110110110001111" when sig_inp <= "000000000000000000000001001111101001" else
--"0110110100010011" when sig_inp <= "000000000000000000000001010001111010" else
--"0110110010010111" when sig_inp <= "000000000000000000000001010100001100" else
--"0110110000011011" when sig_inp <= "000000000000000000000001010110011110" else
--"0110101110100001" when sig_inp <= "000000000000000000000001011000101111" else
--"0110101100100111" when sig_inp <= "000000000000000000000001011011000001" else
--"0110101010101101" when sig_inp <= "000000000000000000000001011101010011" else
--"0110101000110100" when sig_inp <= "000000000000000000000001011111100100" else
--"0110100110111011" when sig_inp <= "000000000000000000000001100001110110" else
--"0110100101000011" when sig_inp <= "000000000000000000000001100100000111" else
--"0110100011001100" when sig_inp <= "000000000000000000000001100110011001" else
--"0110100001010101" when sig_inp <= "000000000000000000000001101000101011" else
--"0110011111011110" when sig_inp <= "000000000000000000000001101010111100" else
--"0110011101101000" when sig_inp <= "000000000000000000000001101101001110" else
--"0110011011110011" when sig_inp <= "000000000000000000000001101111100000" else
--"0110011001111110" when sig_inp <= "000000000000000000000001110001110001" else
--"0110011000001010" when sig_inp <= "000000000000000000000001110100000011" else
--"0110010110010110" when sig_inp <= "000000000000000000000001110110010101" else
--"0110010100100011" when sig_inp <= "000000000000000000000001111000100110" else
--"0110010010110000" when sig_inp <= "000000000000000000000001111010111000" else
--"0110010000111101" when sig_inp <= "000000000000000000000001111101001001" else
--"0110001111001100" when sig_inp <= "000000000000000000000001111111011011" else
--"0110001101011010" when sig_inp <= "000000000000000000000010000001101101" else
--"0110001011101010" when sig_inp <= "000000000000000000000010000011111110" else
--"0110001001111001" when sig_inp <= "000000000000000000000010000110010000" else
--"0110001000001001" when sig_inp <= "000000000000000000000010001000100010" else
--"0110000110011010" when sig_inp <= "000000000000000000000010001010110011" else
--"0110000100101011" when sig_inp <= "000000000000000000000010001101000101" else
--"0110000010111101" when sig_inp <= "000000000000000000000010001111010111" else
--"0110000001001111" when sig_inp <= "000000000000000000000010010001101000" else
--"0101111111100010" when sig_inp <= "000000000000000000000010010011111010" else
--"0101111101110101" when sig_inp <= "000000000000000000000010010110001011" else
--"0101111100001001" when sig_inp <= "000000000000000000000010011000011101" else
--"0101111010011101" when sig_inp <= "000000000000000000000010011010101111" else
--"0101111000110001" when sig_inp <= "000000000000000000000010011101000000" else
--"0101110111000110" when sig_inp <= "000000000000000000000010011111010010" else
--"0101110101011100" when sig_inp <= "000000000000000000000010100001100100" else
--"0101110011110010" when sig_inp <= "000000000000000000000010100011110101" else
--"0101110010001000" when sig_inp <= "000000000000000000000010100110000111" else
--"0101110000011111" when sig_inp <= "000000000000000000000010101000011001" else
--"0101101110110111" when sig_inp <= "000000000000000000000010101010101010" else
--"0101101101001111" when sig_inp <= "000000000000000000000010101100111100" else
--"0101101011100111" when sig_inp <= "000000000000000000000010101111001101" else
--"0101101010000000" when sig_inp <= "000000000000000000000010110001011111" else
--"0101101000011001" when sig_inp <= "000000000000000000000010110011110001" else
--"0101100110110011" when sig_inp <= "000000000000000000000010110110000010" else
--"0101100101001101" when sig_inp <= "000000000000000000000010111000010100" else
--"0101100011101000" when sig_inp <= "000000000000000000000010111010100110" else
--"0101100010000011" when sig_inp <= "000000000000000000000010111100110111" else
--"0101100000011110" when sig_inp <= "000000000000000000000010111111001001" else
--"0101011110111010" when sig_inp <= "000000000000000000000011000001011011" else
--"0101011101010111" when sig_inp <= "000000000000000000000011000011101100" else
--"0101011011110011" when sig_inp <= "000000000000000000000011000101111110" else
--"0101011010010001" when sig_inp <= "000000000000000000000011001000001111" else
--"0101011000101110" when sig_inp <= "000000000000000000000011001010100001" else
--"0101010111001101" when sig_inp <= "000000000000000000000011001100110011" else
--"0101010101101011" when sig_inp <= "000000000000000000000011001111000100" else
--"0101010100001010" when sig_inp <= "000000000000000000000011010001010110" else
--"0101010010101010" when sig_inp <= "000000000000000000000011010011101000" else
--"0101010001001010" when sig_inp <= "000000000000000000000011010101111001" else
--"0101001111101010" when sig_inp <= "000000000000000000000011011000001011" else
--"0101001110001011" when sig_inp <= "000000000000000000000011011010011101" else
--"0101001100101100" when sig_inp <= "000000000000000000000011011100101110" else
--"0101001011001101" when sig_inp <= "000000000000000000000011011111000000" else
--"0101001001101111" when sig_inp <= "000000000000000000000011100001010001" else
--"0101001000010010" when sig_inp <= "000000000000000000000011100011100011" else
--"0101000110110101" when sig_inp <= "000000000000000000000011100101110101" else
--"0101000101011000" when sig_inp <= "000000000000000000000011101000000110" else
--"0101000011111011" when sig_inp <= "000000000000000000000011101010011000" else
--"0101000010011111" when sig_inp <= "000000000000000000000011101100101010" else
--"0101000001000100" when sig_inp <= "000000000000000000000011101110111011" else
--"0100111111101001" when sig_inp <= "000000000000000000000011110001001101" else
--"0100111110001110" when sig_inp <= "000000000000000000000011110011011111" else
--"0100111100110100" when sig_inp <= "000000000000000000000011110101110000" else
--"0100111011011010" when sig_inp <= "000000000000000000000011111000000010" else
--"0100111010000000" when sig_inp <= "000000000000000000000011111010010011" else
--"0100111000100111" when sig_inp <= "000000000000000000000011111100100101" else
--"0100110111001111" when sig_inp <= "000000000000000000000011111110110111" else
--"0100110101110110" when sig_inp <= "000000000000000000000100000001001000" else
--"0100110100011110" when sig_inp <= "000000000000000000000100000011011010" else
--"0100110011000111" when sig_inp <= "000000000000000000000100000101101100" else
--"0100110001110000" when sig_inp <= "000000000000000000000100000111111101" else
--"0100110000011001" when sig_inp <= "000000000000000000000100001010001111" else
--"0100101111000010" when sig_inp <= "000000000000000000000100001100100000" else
--"0100101101101100" when sig_inp <= "000000000000000000000100001110110010" else
--"0100101100010111" when sig_inp <= "000000000000000000000100010001000100" else
--"0100101011000001" when sig_inp <= "000000000000000000000100010011010101" else
--"0100101001101101" when sig_inp <= "000000000000000000000100010101100111" else
--"0100101000011000" when sig_inp <= "000000000000000000000100010111111001" else
--"0100100111000100" when sig_inp <= "000000000000000000000100011010001010" else
--"0100100101110000" when sig_inp <= "000000000000000000000100011100011100" else
--"0100100100011101" when sig_inp <= "000000000000000000000100011110101110" else
--"0100100011001010" when sig_inp <= "000000000000000000000100100000111111" else
--"0100100001110111" when sig_inp <= "000000000000000000000100100011010001" else
--"0100100000100101" when sig_inp <= "000000000000000000000100100101100010" else
--"0100011111010011" when sig_inp <= "000000000000000000000100100111110100" else
--"0100011110000010" when sig_inp <= "000000000000000000000100101010000110" else
--"0100011100110000" when sig_inp <= "000000000000000000000100101100010111" else
--"0100011011100000" when sig_inp <= "000000000000000000000100101110101001" else
--"0100011010001111" when sig_inp <= "000000000000000000000100110000111011" else
--"0100011000111111" when sig_inp <= "000000000000000000000100110011001100" else
--"0100010111101111" when sig_inp <= "000000000000000000000100110101011110" else
--"0100010110100000" when sig_inp <= "000000000000000000000100110111110000" else
--"0100010101010001" when sig_inp <= "000000000000000000000100111010000001" else
--"0100010100000010" when sig_inp <= "000000000000000000000100111100010011" else
--"0100010010110100" when sig_inp <= "000000000000000000000100111110100100" else
--"0100010001100110" when sig_inp <= "000000000000000000000101000000110110" else
--"0100010000011000" when sig_inp <= "000000000000000000000101000011001000" else
--"0100001111001011" when sig_inp <= "000000000000000000000101000101011001" else
--"0100001101111110" when sig_inp <= "000000000000000000000101000111101011" else
--"0100001100110001" when sig_inp <= "000000000000000000000101001001111101" else
--"0100001011100101" when sig_inp <= "000000000000000000000101001100001110" else
--"0100001010011001" when sig_inp <= "000000000000000000000101001110100000" else
--"0100001001001101" when sig_inp <= "000000000000000000000101010000110010" else
--"0100001000000010" when sig_inp <= "000000000000000000000101010011000011" else
--"0100000110110111" when sig_inp <= "000000000000000000000101010101010101" else
--"0100000101101101" when sig_inp <= "000000000000000000000101010111100110" else
--"0100000100100010" when sig_inp <= "000000000000000000000101011001111000" else
--"0100000011011000" when sig_inp <= "000000000000000000000101011100001010" else
--"0100000010001111" when sig_inp <= "000000000000000000000101011110011011" else
--"0100000001000101" when sig_inp <= "000000000000000000000101100000101101" else
--"0011111111111100" when sig_inp <= "000000000000000000000101100010111111" else
--"0011111110110100" when sig_inp <= "000000000000000000000101100101010000" else
--"0011111101101011" when sig_inp <= "000000000000000000000101100111100010" else
--"0011111100100011" when sig_inp <= "000000000000000000000101101001110100" else
--"0011111011011100" when sig_inp <= "000000000000000000000101101100000101" else
--"0011111010010100" when sig_inp <= "000000000000000000000101101110010111" else
--"0011111001001101" when sig_inp <= "000000000000000000000101110000101000" else
--"0011111000000111" when sig_inp <= "000000000000000000000101110010111010" else
--"0011110111000000" when sig_inp <= "000000000000000000000101110101001100" else
--"0011110101111010" when sig_inp <= "000000000000000000000101110111011101" else
--"0011110100110100" when sig_inp <= "000000000000000000000101111001101111" else
--"0011110011101111" when sig_inp <= "000000000000000000000101111100000001" else
--"0011110010101010" when sig_inp <= "000000000000000000000101111110010010" else
--"0011110001100101" when sig_inp <= "000000000000000000000110000000100100" else
--"0011110000100000" when sig_inp <= "000000000000000000000110000010110110" else
--"0011101111011100" when sig_inp <= "000000000000000000000110000101000111" else
--"0011101110011000" when sig_inp <= "000000000000000000000110000111011001" else
--"0011101101010100" when sig_inp <= "000000000000000000000110001001101010" else
--"0011101100010001" when sig_inp <= "000000000000000000000110001011111100" else
--"0011101011001110" when sig_inp <= "000000000000000000000110001110001110" else
--"0011101010001011" when sig_inp <= "000000000000000000000110010000011111" else
--"0011101001001001" when sig_inp <= "000000000000000000000110010010110001" else
--"0011101000000111" when sig_inp <= "000000000000000000000110010101000011" else
--"0011100111000101" when sig_inp <= "000000000000000000000110010111010100" else
--"0011100110000011" when sig_inp <= "000000000000000000000110011001100110" else
--"0011100101000010" when sig_inp <= "000000000000000000000110011011111000" else
--"0011100100000001" when sig_inp <= "000000000000000000000110011110001001" else
--"0011100011000000" when sig_inp <= "000000000000000000000110100000011011" else
--"0011100010000000" when sig_inp <= "000000000000000000000110100010101100" else
--"0011100001000000" when sig_inp <= "000000000000000000000110100100111110" else
--"0011100000000000" when sig_inp <= "000000000000000000000110100111010000" else
--"0011011111000000" when sig_inp <= "000000000000000000000110101001100001" else
--"0011011110000001" when sig_inp <= "000000000000000000000110101011110011" else
--"0011011101000010" when sig_inp <= "000000000000000000000110101110000101" else
--"0011011100000011" when sig_inp <= "000000000000000000000110110000010110" else
--"0011011011000101" when sig_inp <= "000000000000000000000110110010101000" else
--"0011011010000110" when sig_inp <= "000000000000000000000110110100111010" else
--"0011011001001001" when sig_inp <= "000000000000000000000110110111001011" else
--"0011011000001011" when sig_inp <= "000000000000000000000110111001011101" else
--"0011010111001110" when sig_inp <= "000000000000000000000110111011101110" else
--"0011010110010000" when sig_inp <= "000000000000000000000110111110000000" else
--"0011010101010100" when sig_inp <= "000000000000000000000111000000010010" else
--"0011010100010111" when sig_inp <= "000000000000000000000111000010100011" else
--"0011010011011011" when sig_inp <= "000000000000000000000111000100110101" else
--"0011010010011111" when sig_inp <= "000000000000000000000111000111000111" else
--"0011010001100011" when sig_inp <= "000000000000000000000111001001011000" else
--"0011010000101000" when sig_inp <= "000000000000000000000111001011101010" else
--"0011001111101100" when sig_inp <= "000000000000000000000111001101111100" else
--"0011001110110001" when sig_inp <= "000000000000000000000111010000001101" else
--"0011001101110111" when sig_inp <= "000000000000000000000111010010011111" else
--"0011001100111100" when sig_inp <= "000000000000000000000111010100110000" else
--"0011001100000010" when sig_inp <= "000000000000000000000111010111000010" else
--"0011001011001000" when sig_inp <= "000000000000000000000111011001010100" else
--"0011001010001111" when sig_inp <= "000000000000000000000111011011100101" else
--"0011001001010101" when sig_inp <= "000000000000000000000111011101110111" else
--"0011001000011100" when sig_inp <= "000000000000000000000111100000001001" else
--"0011000111100011" when sig_inp <= "000000000000000000000111100010011010" else
--"0011000110101011" when sig_inp <= "000000000000000000000111100100101100" else
--"0011000101110010" when sig_inp <= "000000000000000000000111100110111110" else
--"0011000100111010" when sig_inp <= "000000000000000000000111101001001111" else
--"0011000100000010" when sig_inp <= "000000000000000000000111101011100001" else
--"0011000011001010" when sig_inp <= "000000000000000000000111101101110010" else
--"0011000010010011" when sig_inp <= "000000000000000000000111110000000100" else
--"0011000001011100" when sig_inp <= "000000000000000000000111110010010110" else
--"0011000000100101" when sig_inp <= "000000000000000000000111110100100111" else
--"0010111111101110" when sig_inp <= "000000000000000000000111110110111001" else
--"0010111110111000" when sig_inp <= "000000000000000000000111111001001011" else
--"0010111110000010" when sig_inp <= "000000000000000000000111111011011100" else
--"0010111101001100" when sig_inp <= "000000000000000000000111111101101110" else
--"0010111100010110" when sig_inp <= "000000000000000000001000000000000000" else
--"0010111011100001" when sig_inp <= "000000000000000000001000000010010001" else
--"0010111010101011" when sig_inp <= "000000000000000000001000000100100011" else
--"0010111001110111" when sig_inp <= "000000000000000000001000000110110100" else
--"0010111001000010" when sig_inp <= "000000000000000000001000001001000110" else
--"0010111000001101" when sig_inp <= "000000000000000000001000001011011000" else
--"0010110111011001" when sig_inp <= "000000000000000000001000001101101001" else
--"0010110110100101" when sig_inp <= "000000000000000000001000001111111011" else
--"0010110101110001" when sig_inp <= "000000000000000000001000010010001101" else
--"0010110100111110" when sig_inp <= "000000000000000000001000010100011110" else
--"0010110100001010" when sig_inp <= "000000000000000000001000010110110000" else
--"0010110011010111" when sig_inp <= "000000000000000000001000011001000001" else
--"0010110010100100" when sig_inp <= "000000000000000000001000011011010011" else
--"0010110001110001" when sig_inp <= "000000000000000000001000011101100101" else
--"0010110000111111" when sig_inp <= "000000000000000000001000011111110110" else
--"0010110000001101" when sig_inp <= "000000000000000000001000100010001000" else
--"0010101111011011" when sig_inp <= "000000000000000000001000100100011010" else
--"0010101110101001" when sig_inp <= "000000000000000000001000100110101011" else
--"0010101101110111" when sig_inp <= "000000000000000000001000101000111101" else
--"0010101101000110" when sig_inp <= "000000000000000000001000101011001111" else
--"0010101100010101" when sig_inp <= "000000000000000000001000101101100000" else
--"0010101011100100" when sig_inp <= "000000000000000000001000101111110010" else
--"0010101010110011" when sig_inp <= "000000000000000000001000110010000011" else
--"0010101010000011" when sig_inp <= "000000000000000000001000110100010101" else
--"0010101001010011" when sig_inp <= "000000000000000000001000110110100111" else
--"0010101000100010" when sig_inp <= "000000000000000000001000111000111000" else
--"0010100111110011" when sig_inp <= "000000000000000000001000111011001010" else
--"0010100111000011" when sig_inp <= "000000000000000000001000111101011100" else
--"0010100110010100" when sig_inp <= "000000000000000000001000111111101101" else
--"0010100101100100" when sig_inp <= "000000000000000000001001000001111111" else
--"0010100100110101" when sig_inp <= "000000000000000000001001000100010001" else
--"0010100100000111" when sig_inp <= "000000000000000000001001000110100010" else
--"0010100011011000" when sig_inp <= "000000000000000000001001001000110100" else
--"0010100010101010" when sig_inp <= "000000000000000000001001001011000101" else
--"0010100001111100" when sig_inp <= "000000000000000000001001001101010111" else
--"0010100001001110" when sig_inp <= "000000000000000000001001001111101001" else
--"0010100000100000" when sig_inp <= "000000000000000000001001010001111010" else
--"0010011111110010" when sig_inp <= "000000000000000000001001010100001100" else
--"0010011111000101" when sig_inp <= "000000000000000000001001010110011110" else
--"0010011110011000" when sig_inp <= "000000000000000000001001011000101111" else
--"0010011101101011" when sig_inp <= "000000000000000000001001011011000001" else
--"0010011100111110" when sig_inp <= "000000000000000000001001011101010011" else
--"0010011100010010" when sig_inp <= "000000000000000000001001011111100100" else
--"0010011011100101" when sig_inp <= "000000000000000000001001100001110110" else
--"0010011010111001" when sig_inp <= "000000000000000000001001100100000111" else
--"0010011010001101" when sig_inp <= "000000000000000000001001100110011001" else
--"0010011001100001" when sig_inp <= "000000000000000000001001101000101011" else
--"0010011000110110" when sig_inp <= "000000000000000000001001101010111100" else
--"0010011000001010" when sig_inp <= "000000000000000000001001101101001110" else
--"0010010111011111" when sig_inp <= "000000000000000000001001101111100000" else
--"0010010110110100" when sig_inp <= "000000000000000000001001110001110001" else
--"0010010110001001" when sig_inp <= "000000000000000000001001110100000011" else
--"0010010101011111" when sig_inp <= "000000000000000000001001110110010101" else
--"0010010100110100" when sig_inp <= "000000000000000000001001111000100110" else
--"0010010100001010" when sig_inp <= "000000000000000000001001111010111000" else
--"0010010011100000" when sig_inp <= "000000000000000000001001111101001001" else
--"0010010010110110" when sig_inp <= "000000000000000000001001111111011011" else
--"0010010010001100" when sig_inp <= "000000000000000000001010000001101101" else
--"0010010001100011" when sig_inp <= "000000000000000000001010000011111110" else
--"0010010000111010" when sig_inp <= "000000000000000000001010000110010000" else
--"0010010000010001" when sig_inp <= "000000000000000000001010001000100010" else
--"0010001111101000" when sig_inp <= "000000000000000000001010001010110011" else
--"0010001110111111" when sig_inp <= "000000000000000000001010001101000101" else
--"0010001110010110" when sig_inp <= "000000000000000000001010001111010111" else
--"0010001101101110" when sig_inp <= "000000000000000000001010010001101000" else
--"0010001101000110" when sig_inp <= "000000000000000000001010010011111010" else
--"0010001100011110" when sig_inp <= "000000000000000000001010010110001011" else
--"0010001011110110" when sig_inp <= "000000000000000000001010011000011101" else
--"0010001011001110" when sig_inp <= "000000000000000000001010011010101111" else
--"0010001010100110" when sig_inp <= "000000000000000000001010011101000000" else
--"0010001001111111" when sig_inp <= "000000000000000000001010011111010010" else
--"0010001001011000" when sig_inp <= "000000000000000000001010100001100100" else
--"0010001000110001" when sig_inp <= "000000000000000000001010100011110101" else
--"0010001000001010" when sig_inp <= "000000000000000000001010100110000111" else
--"0010000111100100" when sig_inp <= "000000000000000000001010101000011001" else
--"0010000110111101" when sig_inp <= "000000000000000000001010101010101010" else
--"0010000110010111" when sig_inp <= "000000000000000000001010101100111100" else
--"0010000101110001" when sig_inp <= "000000000000000000001010101111001101" else
--"0010000101001011" when sig_inp <= "000000000000000000001010110001011111" else
--"0010000100100101" when sig_inp <= "000000000000000000001010110011110001" else
--"0010000011111111" when sig_inp <= "000000000000000000001010110110000010" else
--"0010000011011010" when sig_inp <= "000000000000000000001010111000010100" else
--"0010000010110100" when sig_inp <= "000000000000000000001010111010100110" else
--"0010000010001111" when sig_inp <= "000000000000000000001010111100110111" else
--"0010000001101010" when sig_inp <= "000000000000000000001010111111001001" else
--"0010000001000110" when sig_inp <= "000000000000000000001011000001011011" else
--"0010000000100001" when sig_inp <= "000000000000000000001011000011101100" else
--"0001111111111100" when sig_inp <= "000000000000000000001011000101111110" else
--"0001111111011000" when sig_inp <= "000000000000000000001011001000001111" else
--"0001111110110100" when sig_inp <= "000000000000000000001011001010100001" else
--"0001111110010000" when sig_inp <= "000000000000000000001011001100110011" else
--"0001111101101100" when sig_inp <= "000000000000000000001011001111000100" else
--"0001111101001000" when sig_inp <= "000000000000000000001011010001010110" else
--"0001111100100101" when sig_inp <= "000000000000000000001011010011101000" else
--"0001111100000010" when sig_inp <= "000000000000000000001011010101111001" else
--"0001111011011110" when sig_inp <= "000000000000000000001011011000001011" else
--"0001111010111011" when sig_inp <= "000000000000000000001011011010011101" else
--"0001111010011000" when sig_inp <= "000000000000000000001011011100101110" else
--"0001111001110110" when sig_inp <= "000000000000000000001011011111000000" else
--"0001111001010011" when sig_inp <= "000000000000000000001011100001010001" else
--"0001111000110001" when sig_inp <= "000000000000000000001011100011100011" else
--"0001111000001110" when sig_inp <= "000000000000000000001011100101110101" else
--"0001110111101100" when sig_inp <= "000000000000000000001011101000000110" else
--"0001110111001010" when sig_inp <= "000000000000000000001011101010011000" else
--"0001110110101001" when sig_inp <= "000000000000000000001011101100101010" else
--"0001110110000111" when sig_inp <= "000000000000000000001011101110111011" else
--"0001110101100101" when sig_inp <= "000000000000000000001011110001001101" else
--"0001110101000100" when sig_inp <= "000000000000000000001011110011011111" else
--"0001110100100011" when sig_inp <= "000000000000000000001011110101110000" else
--"0001110100000010" when sig_inp <= "000000000000000000001011111000000010" else
--"0001110011100001" when sig_inp <= "000000000000000000001011111010010011" else
--"0001110011000000" when sig_inp <= "000000000000000000001011111100100101" else
--"0001110010011111" when sig_inp <= "000000000000000000001011111110110111" else
--"0001110001111111" when sig_inp <= "000000000000000000001100000001001000" else
--"0001110001011110" when sig_inp <= "000000000000000000001100000011011010" else
--"0001110000111110" when sig_inp <= "000000000000000000001100000101101100" else
--"0001110000011110" when sig_inp <= "000000000000000000001100000111111101" else
--"0001101111111110" when sig_inp <= "000000000000000000001100001010001111" else
--"0001101111011110" when sig_inp <= "000000000000000000001100001100100000" else
--"0001101110111111" when sig_inp <= "000000000000000000001100001110110010" else
--"0001101110011111" when sig_inp <= "000000000000000000001100010001000100" else
--"0001101110000000" when sig_inp <= "000000000000000000001100010011010101" else
--"0001101101100001" when sig_inp <= "000000000000000000001100010101100111" else
--"0001101101000010" when sig_inp <= "000000000000000000001100010111111001" else
--"0001101100100011" when sig_inp <= "000000000000000000001100011010001010" else
--"0001101100000100" when sig_inp <= "000000000000000000001100011100011100" else
--"0001101011100101" when sig_inp <= "000000000000000000001100011110101110" else
--"0001101011000111" when sig_inp <= "000000000000000000001100100000111111" else
--"0001101010101000" when sig_inp <= "000000000000000000001100100011010001" else
--"0001101010001010" when sig_inp <= "000000000000000000001100100101100010" else
--"0001101001101100" when sig_inp <= "000000000000000000001100100111110100" else
--"0001101001001110" when sig_inp <= "000000000000000000001100101010000110" else
--"0001101000110000" when sig_inp <= "000000000000000000001100101100010111" else
--"0001101000010010" when sig_inp <= "000000000000000000001100101110101001" else
--"0001100111110101" when sig_inp <= "000000000000000000001100110000111011" else
--"0001100111010111" when sig_inp <= "000000000000000000001100110011001100" else
--"0001100110111010" when sig_inp <= "000000000000000000001100110101011110" else
--"0001100110011101" when sig_inp <= "000000000000000000001100110111110000" else
--"0001100110000000" when sig_inp <= "000000000000000000001100111010000001" else
--"0001100101100011" when sig_inp <= "000000000000000000001100111100010011" else
--"0001100101000110" when sig_inp <= "000000000000000000001100111110100100" else
--"0001100100101001" when sig_inp <= "000000000000000000001101000000110110" else
--"0001100100001101" when sig_inp <= "000000000000000000001101000011001000" else
--"0001100011110000" when sig_inp <= "000000000000000000001101000101011001" else
--"0001100011010100" when sig_inp <= "000000000000000000001101000111101011" else
--"0001100010111000" when sig_inp <= "000000000000000000001101001001111101" else
--"0001100010011100" when sig_inp <= "000000000000000000001101001100001110" else
--"0001100010000000" when sig_inp <= "000000000000000000001101001110100000" else
--"0001100001100100" when sig_inp <= "000000000000000000001101010000110010" else
--"0001100001001000" when sig_inp <= "000000000000000000001101010011000011" else
--"0001100000101101" when sig_inp <= "000000000000000000001101010101010101" else
--"0001100000010001" when sig_inp <= "000000000000000000001101010111100110" else
--"0001011111110110" when sig_inp <= "000000000000000000001101011001111000" else
--"0001011111011011" when sig_inp <= "000000000000000000001101011100001010" else
--"0001011111000000" when sig_inp <= "000000000000000000001101011110011011" else
--"0001011110100101" when sig_inp <= "000000000000000000001101100000101101" else
--"0001011110001010" when sig_inp <= "000000000000000000001101100010111111" else
--"0001011101101111" when sig_inp <= "000000000000000000001101100101010000" else
--"0001011101010100" when sig_inp <= "000000000000000000001101100111100010" else
--"0001011100111010" when sig_inp <= "000000000000000000001101101001110100" else
--"0001011100100000" when sig_inp <= "000000000000000000001101101100000101" else
--"0001011100000101" when sig_inp <= "000000000000000000001101101110010111" else
--"0001011011101011" when sig_inp <= "000000000000000000001101110000101000" else
--"0001011011010001" when sig_inp <= "000000000000000000001101110010111010" else
--"0001011010110111" when sig_inp <= "000000000000000000001101110101001100" else
--"0001011010011101" when sig_inp <= "000000000000000000001101110111011101" else
--"0001011010000100" when sig_inp <= "000000000000000000001101111001101111" else
--"0001011001101010" when sig_inp <= "000000000000000000001101111100000001" else
--"0001011001010001" when sig_inp <= "000000000000000000001101111110010010" else
--"0001011000110111" when sig_inp <= "000000000000000000001110000000100100" else
--"0001011000011110" when sig_inp <= "000000000000000000001110000010110110" else
--"0001011000000101" when sig_inp <= "000000000000000000001110000101000111" else
--"0001010111101100" when sig_inp <= "000000000000000000001110000111011001" else
--"0001010111010011" when sig_inp <= "000000000000000000001110001001101010" else
--"0001010110111010" when sig_inp <= "000000000000000000001110001011111100" else
--"0001010110100010" when sig_inp <= "000000000000000000001110001110001110" else
--"0001010110001001" when sig_inp <= "000000000000000000001110010000011111" else
--"0001010101110001" when sig_inp <= "000000000000000000001110010010110001" else
--"0001010101011000" when sig_inp <= "000000000000000000001110010101000011" else
--"0001010101000000" when sig_inp <= "000000000000000000001110010111010100" else
--"0001010100101000" when sig_inp <= "000000000000000000001110011001100110" else
--"0001010100010000" when sig_inp <= "000000000000000000001110011011111000" else
--"0001010011111000" when sig_inp <= "000000000000000000001110011110001001" else
--"0001010011100000" when sig_inp <= "000000000000000000001110100000011011" else
--"0001010011001001" when sig_inp <= "000000000000000000001110100010101100" else
--"0001010010110001" when sig_inp <= "000000000000000000001110100100111110" else
--"0001010010011001" when sig_inp <= "000000000000000000001110100111010000" else
--"0001010010000010" when sig_inp <= "000000000000000000001110101001100001" else
--"0001010001101011" when sig_inp <= "000000000000000000001110101011110011" else
--"0001010001010100" when sig_inp <= "000000000000000000001110101110000101" else
--"0001010000111101" when sig_inp <= "000000000000000000001110110000010110" else
--"0001010000100110" when sig_inp <= "000000000000000000001110110010101000" else
--"0001010000001111" when sig_inp <= "000000000000000000001110110100111010" else
--"0001001111111000" when sig_inp <= "000000000000000000001110110111001011" else
--"0001001111100001" when sig_inp <= "000000000000000000001110111001011101" else
--"0001001111001011" when sig_inp <= "000000000000000000001110111011101110" else
--"0001001110110100" when sig_inp <= "000000000000000000001110111110000000" else
--"0001001110011110" when sig_inp <= "000000000000000000001111000000010010" else
--"0001001110001000" when sig_inp <= "000000000000000000001111000010100011" else
--"0001001101110001" when sig_inp <= "000000000000000000001111000100110101" else
--"0001001101011011" when sig_inp <= "000000000000000000001111000111000111" else
--"0001001101000101" when sig_inp <= "000000000000000000001111001001011000" else
--"0001001100101111" when sig_inp <= "000000000000000000001111001011101010" else
--"0001001100011010" when sig_inp <= "000000000000000000001111001101111100" else
--"0001001100000100" when sig_inp <= "000000000000000000001111010000001101" else
--"0001001011101110" when sig_inp <= "000000000000000000001111010010011111" else
--"0001001011011001" when sig_inp <= "000000000000000000001111010100110000" else
--"0001001011000100" when sig_inp <= "000000000000000000001111010111000010" else
--"0001001010101110" when sig_inp <= "000000000000000000001111011001010100" else
--"0001001010011001" when sig_inp <= "000000000000000000001111011011100101" else
--"0001001010000100" when sig_inp <= "000000000000000000001111011101110111" else
--"0001001001101111" when sig_inp <= "000000000000000000001111100000001001" else
--"0001001001011010" when sig_inp <= "000000000000000000001111100010011010" else
--"0001001001000101" when sig_inp <= "000000000000000000001111100100101100" else
--"0001001000110000" when sig_inp <= "000000000000000000001111100110111110" else
--"0001001000011100" when sig_inp <= "000000000000000000001111101001001111" else
--"0001001000000111" when sig_inp <= "000000000000000000001111101011100001" else
--"0001000111110011" when sig_inp <= "000000000000000000001111101101110010" else
--"0001000111011110" when sig_inp <= "000000000000000000001111110000000100" else
--"0001000111001010" when sig_inp <= "000000000000000000001111110010010110" else
--"0001000110110110" when sig_inp <= "000000000000000000001111110100100111" else
--"0001000110100010" when sig_inp <= "000000000000000000001111110110111001" else
--"0001000110001110" when sig_inp <= "000000000000000000001111111001001011" else
--"0001000101111010" when sig_inp <= "000000000000000000001111111011011100" else
--"0001000101100110" when sig_inp <= "000000000000000000001111111101101110" else
--"0001000101010010" when sig_inp <= "000000000000000000010000000000000000" else
--"0001000100111111" when sig_inp <= "000000000000000000010000000010010001" else
--"0001000100101011" when sig_inp <= "000000000000000000010000000100100011" else
--"0001000100010111" when sig_inp <= "000000000000000000010000000110110100" else
--"0001000100000100" when sig_inp <= "000000000000000000010000001001000110" else
--"0001000011110001" when sig_inp <= "000000000000000000010000001011011000" else
--"0001000011011101" when sig_inp <= "000000000000000000010000001101101001" else
--"0001000011001010" when sig_inp <= "000000000000000000010000001111111011" else
--"0001000010110111" when sig_inp <= "000000000000000000010000010010001101" else
--"0001000010100100" when sig_inp <= "000000000000000000010000010100011110" else
--"0001000010010001" when sig_inp <= "000000000000000000010000010110110000" else
--"0001000001111111" when sig_inp <= "000000000000000000010000011001000001" else
--"0001000001101100" when sig_inp <= "000000000000000000010000011011010011" else
--"0001000001011001" when sig_inp <= "000000000000000000010000011101100101" else
--"0001000001000111" when sig_inp <= "000000000000000000010000011111110110" else
--"0001000000110100" when sig_inp <= "000000000000000000010000100010001000" else
--"0001000000100010" when sig_inp <= "000000000000000000010000100100011010" else
--"0001000000001111" when sig_inp <= "000000000000000000010000100110101011" else
--"0000111111111101" when sig_inp <= "000000000000000000010000101000111101" else
--"0000111111101011" when sig_inp <= "000000000000000000010000101011001111" else
--"0000111111011001" when sig_inp <= "000000000000000000010000101101100000" else
--"0000111111000111" when sig_inp <= "000000000000000000010000101111110010" else
--"0000111110110101" when sig_inp <= "000000000000000000010000110010000011" else
--"0000111110100011" when sig_inp <= "000000000000000000010000110100010101" else
--"0000111110010001" when sig_inp <= "000000000000000000010000110110100111" else
--"0000111110000000" when sig_inp <= "000000000000000000010000111000111000" else
--"0000111101101110" when sig_inp <= "000000000000000000010000111011001010" else
--"0000111101011101" when sig_inp <= "000000000000000000010000111101011100" else
--"0000111101001011" when sig_inp <= "000000000000000000010000111111101101" else
--"0000111100111010" when sig_inp <= "000000000000000000010001000001111111" else
--"0000111100101001" when sig_inp <= "000000000000000000010001000100010001" else
--"0000111100010111" when sig_inp <= "000000000000000000010001000110100010" else
--"0000111100000110" when sig_inp <= "000000000000000000010001001000110100" else
--"0000111011110101" when sig_inp <= "000000000000000000010001001011000101" else
--"0000111011100100" when sig_inp <= "000000000000000000010001001101010111" else
--"0000111011010011" when sig_inp <= "000000000000000000010001001111101001" else
--"0000111011000010" when sig_inp <= "000000000000000000010001010001111010" else
--"0000111010110010" when sig_inp <= "000000000000000000010001010100001100" else
--"0000111010100001" when sig_inp <= "000000000000000000010001010110011110" else
--"0000111010010000" when sig_inp <= "000000000000000000010001011000101111" else
--"0000111010000000" when sig_inp <= "000000000000000000010001011011000001" else
--"0000111001101111" when sig_inp <= "000000000000000000010001011101010011" else
--"0000111001011111" when sig_inp <= "000000000000000000010001011111100100" else
--"0000111001001111" when sig_inp <= "000000000000000000010001100001110110" else
--"0000111000111110" when sig_inp <= "000000000000000000010001100100000111" else
--"0000111000101110" when sig_inp <= "000000000000000000010001100110011001" else
--"0000111000011110" when sig_inp <= "000000000000000000010001101000101011" else
--"0000111000001110" when sig_inp <= "000000000000000000010001101010111100" else
--"0000110111111110" when sig_inp <= "000000000000000000010001101101001110" else
--"0000110111101110" when sig_inp <= "000000000000000000010001101111100000" else
--"0000110111011111" when sig_inp <= "000000000000000000010001110001110001" else
--"0000110111001111" when sig_inp <= "000000000000000000010001110100000011" else
--"0000110110111111" when sig_inp <= "000000000000000000010001110110010101" else
--"0000110110101111" when sig_inp <= "000000000000000000010001111000100110" else
--"0000110110100000" when sig_inp <= "000000000000000000010001111010111000" else
--"0000110110010000" when sig_inp <= "000000000000000000010001111101001001" else
--"0000110110000001" when sig_inp <= "000000000000000000010001111111011011" else
--"0000110101110010" when sig_inp <= "000000000000000000010010000001101101" else
--"0000110101100010" when sig_inp <= "000000000000000000010010000011111110" else
--"0000110101010011" when sig_inp <= "000000000000000000010010000110010000" else
--"0000110101000100" when sig_inp <= "000000000000000000010010001000100010" else
--"0000110100110101" when sig_inp <= "000000000000000000010010001010110011" else
--"0000110100100110" when sig_inp <= "000000000000000000010010001101000101" else
--"0000110100010111" when sig_inp <= "000000000000000000010010001111010111" else
--"0000110100001000" when sig_inp <= "000000000000000000010010010001101000" else
--"0000110011111001" when sig_inp <= "000000000000000000010010010011111010" else
--"0000110011101011" when sig_inp <= "000000000000000000010010010110001011" else
--"0000110011011100" when sig_inp <= "000000000000000000010010011000011101" else
--"0000110011001101" when sig_inp <= "000000000000000000010010011010101111" else
--"0000110010111111" when sig_inp <= "000000000000000000010010011101000000" else
--"0000110010110000" when sig_inp <= "000000000000000000010010011111010010" else
--"0000110010100010" when sig_inp <= "000000000000000000010010100001100100" else
--"0000110010010100" when sig_inp <= "000000000000000000010010100011110101" else
--"0000110010000101" when sig_inp <= "000000000000000000010010100110000111" else
--"0000110001110111" when sig_inp <= "000000000000000000010010101000011001" else
--"0000110001101001" when sig_inp <= "000000000000000000010010101010101010" else
--"0000110001011011" when sig_inp <= "000000000000000000010010101100111100" else
--"0000110001001101" when sig_inp <= "000000000000000000010010101111001101" else
--"0000110000111111" when sig_inp <= "000000000000000000010010110001011111" else
--"0000110000110001" when sig_inp <= "000000000000000000010010110011110001" else
--"0000110000100011" when sig_inp <= "000000000000000000010010110110000010" else
--"0000110000010101" when sig_inp <= "000000000000000000010010111000010100" else
--"0000110000001000" when sig_inp <= "000000000000000000010010111010100110" else
--"0000101111111010" when sig_inp <= "000000000000000000010010111100110111" else
--"0000101111101100" when sig_inp <= "000000000000000000010010111111001001" else
--"0000101111011111" when sig_inp <= "000000000000000000010011000001011011" else
--"0000101111010001" when sig_inp <= "000000000000000000010011000011101100" else
--"0000101111000100" when sig_inp <= "000000000000000000010011000101111110" else
--"0000101110110111" when sig_inp <= "000000000000000000010011001000001111" else
--"0000101110101001" when sig_inp <= "000000000000000000010011001010100001" else
--"0000101110011100" when sig_inp <= "000000000000000000010011001100110011" else
--"0000101110001111" when sig_inp <= "000000000000000000010011001111000100" else
--"0000101110000010" when sig_inp <= "000000000000000000010011010001010110" else
--"0000101101110101" when sig_inp <= "000000000000000000010011010011101000" else
--"0000101101101000" when sig_inp <= "000000000000000000010011010101111001" else
--"0000101101011011" when sig_inp <= "000000000000000000010011011000001011" else
--"0000101101001110" when sig_inp <= "000000000000000000010011011010011101" else
--"0000101101000001" when sig_inp <= "000000000000000000010011011100101110" else
--"0000101100110100" when sig_inp <= "000000000000000000010011011111000000" else
--"0000101100101000" when sig_inp <= "000000000000000000010011100001010001" else
--"0000101100011011" when sig_inp <= "000000000000000000010011100011100011" else
--"0000101100001110" when sig_inp <= "000000000000000000010011100101110101" else
--"0000101100000010" when sig_inp <= "000000000000000000010011101000000110" else
--"0000101011110101" when sig_inp <= "000000000000000000010011101010011000" else
--"0000101011101001" when sig_inp <= "000000000000000000010011101100101010" else
--"0000101011011100" when sig_inp <= "000000000000000000010011101110111011" else
--"0000101011010000" when sig_inp <= "000000000000000000010011110001001101" else
--"0000101011000100" when sig_inp <= "000000000000000000010011110011011111" else
--"0000101010111000" when sig_inp <= "000000000000000000010011110101110000" else
--"0000101010101011" when sig_inp <= "000000000000000000010011111000000010" else
--"0000101010011111" when sig_inp <= "000000000000000000010011111010010011" else
--"0000101010010011" when sig_inp <= "000000000000000000010011111100100101" else
--"0000101010000111" when sig_inp <= "000000000000000000010011111110110111" else
--"0000101001111011" when sig_inp <= "000000000000000000010100000001001000" else
--"0000101001101111" when sig_inp <= "000000000000000000010100000011011010" else
--"0000101001100100" when sig_inp <= "000000000000000000010100000101101100" else
--"0000101001011000" when sig_inp <= "000000000000000000010100000111111101" else
--"0000101001001100" when sig_inp <= "000000000000000000010100001010001111" else
--"0000101001000000" when sig_inp <= "000000000000000000010100001100100000" else
--"0000101000110101" when sig_inp <= "000000000000000000010100001110110010" else
--"0000101000101001" when sig_inp <= "000000000000000000010100010001000100" else
--"0000101000011110" when sig_inp <= "000000000000000000010100010011010101" else
--"0000101000010010" when sig_inp <= "000000000000000000010100010101100111" else
--"0000101000000111" when sig_inp <= "000000000000000000010100010111111001" else
--"0000100111111011" when sig_inp <= "000000000000000000010100011010001010" else
--"0000100111110000" when sig_inp <= "000000000000000000010100011100011100" else
--"0000100111100101" when sig_inp <= "000000000000000000010100011110101110" else
--"0000100111011001" when sig_inp <= "000000000000000000010100100000111111" else
--"0000100111001110" when sig_inp <= "000000000000000000010100100011010001" else
--"0000100111000011" when sig_inp <= "000000000000000000010100100101100010" else
--"0000100110111000" when sig_inp <= "000000000000000000010100100111110100" else
--"0000100110101101" when sig_inp <= "000000000000000000010100101010000110" else
--"0000100110100010" when sig_inp <= "000000000000000000010100101100010111" else
--"0000100110010111" when sig_inp <= "000000000000000000010100101110101001" else
--"0000100110001100" when sig_inp <= "000000000000000000010100110000111011" else
--"0000100110000001" when sig_inp <= "000000000000000000010100110011001100" else
--"0000100101110111" when sig_inp <= "000000000000000000010100110101011110" else
--"0000100101101100" when sig_inp <= "000000000000000000010100110111110000" else
--"0000100101100001" when sig_inp <= "000000000000000000010100111010000001" else
--"0000100101010110" when sig_inp <= "000000000000000000010100111100010011" else
--"0000100101001100" when sig_inp <= "000000000000000000010100111110100100" else
--"0000100101000001" when sig_inp <= "000000000000000000010101000000110110" else
--"0000100100110111" when sig_inp <= "000000000000000000010101000011001000" else
--"0000100100101100" when sig_inp <= "000000000000000000010101000101011001" else
--"0000100100100010" when sig_inp <= "000000000000000000010101000111101011" else
--"0000100100010111" when sig_inp <= "000000000000000000010101001001111101" else
--"0000100100001101" when sig_inp <= "000000000000000000010101001100001110" else
--"0000100100000011" when sig_inp <= "000000000000000000010101001110100000" else
--"0000100011111001" when sig_inp <= "000000000000000000010101010000110010" else
--"0000100011101110" when sig_inp <= "000000000000000000010101010011000011" else
--"0000100011100100" when sig_inp <= "000000000000000000010101010101010101" else
--"0000100011011010" when sig_inp <= "000000000000000000010101010111100110" else
--"0000100011010000" when sig_inp <= "000000000000000000010101011001111000" else
--"0000100011000110" when sig_inp <= "000000000000000000010101011100001010" else
--"0000100010111100" when sig_inp <= "000000000000000000010101011110011011" else
--"0000100010110010" when sig_inp <= "000000000000000000010101100000101101" else
--"0000100010101000" when sig_inp <= "000000000000000000010101100010111111" else
--"0000100010011111" when sig_inp <= "000000000000000000010101100101010000" else
--"0000100010010101" when sig_inp <= "000000000000000000010101100111100010" else
--"0000100010001011" when sig_inp <= "000000000000000000010101101001110100" else
--"0000100010000001" when sig_inp <= "000000000000000000010101101100000101" else
--"0000100001111000" when sig_inp <= "000000000000000000010101101110010111" else
--"0000100001101110" when sig_inp <= "000000000000000000010101110000101000" else
--"0000100001100101" when sig_inp <= "000000000000000000010101110010111010" else
--"0000100001011011" when sig_inp <= "000000000000000000010101110101001100" else
--"0000100001010001" when sig_inp <= "000000000000000000010101110111011101" else
--"0000100001001000" when sig_inp <= "000000000000000000010101111001101111" else
--"0000100000111111" when sig_inp <= "000000000000000000010101111100000001" else
--"0000100000110101" when sig_inp <= "000000000000000000010101111110010010" else
--"0000100000101100" when sig_inp <= "000000000000000000010110000000100100" else
--"0000100000100011" when sig_inp <= "000000000000000000010110000010110110" else
--"0000100000011001" when sig_inp <= "000000000000000000010110000101000111" else
--"0000100000010000" when sig_inp <= "000000000000000000010110000111011001" else
--"0000100000000111" when sig_inp <= "000000000000000000010110001001101010" else
--"0000011111111110" when sig_inp <= "000000000000000000010110001011111100" else
--"0000011111110101" when sig_inp <= "000000000000000000010110001110001110" else
--"0000011111101100" when sig_inp <= "000000000000000000010110010000011111" else
--"0000011111100011" when sig_inp <= "000000000000000000010110010010110001" else
--"0000011111011010" when sig_inp <= "000000000000000000010110010101000011" else
--"0000011111010001" when sig_inp <= "000000000000000000010110010111010100" else
--"0000011111001000" when sig_inp <= "000000000000000000010110011001100110" else
--"0000011110111111" when sig_inp <= "000000000000000000010110011011111000" else
--"0000011110110110" when sig_inp <= "000000000000000000010110011110001001" else
--"0000011110101110" when sig_inp <= "000000000000000000010110100000011011" else
--"0000011110100101" when sig_inp <= "000000000000000000010110100010101100" else
--"0000011110011100" when sig_inp <= "000000000000000000010110100100111110" else
--"0000011110010100" when sig_inp <= "000000000000000000010110100111010000" else
--"0000011110001011" when sig_inp <= "000000000000000000010110101001100001" else
--"0000011110000011" when sig_inp <= "000000000000000000010110101011110011" else
--"0000011101111010" when sig_inp <= "000000000000000000010110101110000101" else
--"0000011101110010" when sig_inp <= "000000000000000000010110110000010110" else
--"0000011101101001" when sig_inp <= "000000000000000000010110110010101000" else
--"0000011101100001" when sig_inp <= "000000000000000000010110110100111010" else
--"0000011101011000" when sig_inp <= "000000000000000000010110110111001011" else
--"0000011101010000" when sig_inp <= "000000000000000000010110111001011101" else
--"0000011101001000" when sig_inp <= "000000000000000000010110111011101110" else
--"0000011100111111" when sig_inp <= "000000000000000000010110111110000000" else
--"0000011100110111" when sig_inp <= "000000000000000000010111000000010010" else
--"0000011100101111" when sig_inp <= "000000000000000000010111000010100011" else
--"0000011100100111" when sig_inp <= "000000000000000000010111000100110101" else
--"0000011100011111" when sig_inp <= "000000000000000000010111000111000111" else
--"0000011100010111" when sig_inp <= "000000000000000000010111001001011000" else
--"0000011100001111" when sig_inp <= "000000000000000000010111001011101010" else
--"0000011100000110" when sig_inp <= "000000000000000000010111001101111100" else
--"0000011011111111" when sig_inp <= "000000000000000000010111010000001101" else
--"0000011011110111" when sig_inp <= "000000000000000000010111010010011111" else
--"0000011011101111" when sig_inp <= "000000000000000000010111010100110000" else
--"0000011011100111" when sig_inp <= "000000000000000000010111010111000010" else
--"0000011011011111" when sig_inp <= "000000000000000000010111011001010100" else
--"0000011011010111" when sig_inp <= "000000000000000000010111011011100101" else
--"0000011011001111" when sig_inp <= "000000000000000000010111011101110111" else
--"0000011011001000" when sig_inp <= "000000000000000000010111100000001001" else
--"0000011011000000" when sig_inp <= "000000000000000000010111100010011010" else
--"0000011010111000" when sig_inp <= "000000000000000000010111100100101100" else
--"0000011010110001" when sig_inp <= "000000000000000000010111100110111110" else
--"0000011010101001" when sig_inp <= "000000000000000000010111101001001111" else
--"0000011010100010" when sig_inp <= "000000000000000000010111101011100001" else
--"0000011010011010" when sig_inp <= "000000000000000000010111101101110010" else
--"0000011010010010" when sig_inp <= "000000000000000000010111110000000100" else
--"0000011010001011" when sig_inp <= "000000000000000000010111110010010110" else
--"0000011010000100" when sig_inp <= "000000000000000000010111110100100111" else
--"0000011001111100" when sig_inp <= "000000000000000000010111110110111001" else
--"0000011001110101" when sig_inp <= "000000000000000000010111111001001011" else
--"0000011001101101" when sig_inp <= "000000000000000000010111111011011100" else
--"0000011001100110" when sig_inp <= "000000000000000000010111111101101110" else
--"0000011001011111" when sig_inp <= "000000000000000000011000000000000000" else
--"0000011001011000" when sig_inp <= "000000000000000000011000000010010001" else
--"0000011001010000" when sig_inp <= "000000000000000000011000000100100011" else
--"0000011001001001" when sig_inp <= "000000000000000000011000000110110100" else
--"0000011001000010" when sig_inp <= "000000000000000000011000001001000110" else
--"0000011000111011" when sig_inp <= "000000000000000000011000001011011000" else
--"0000011000110100" when sig_inp <= "000000000000000000011000001101101001" else
--"0000011000101101" when sig_inp <= "000000000000000000011000001111111011" else
--"0000011000100110" when sig_inp <= "000000000000000000011000010010001101" else
--"0000011000011111" when sig_inp <= "000000000000000000011000010100011110" else
--"0000011000011000" when sig_inp <= "000000000000000000011000010110110000" else
--"0000011000010001" when sig_inp <= "000000000000000000011000011001000001" else
--"0000011000001010" when sig_inp <= "000000000000000000011000011011010011" else
--"0000011000000011" when sig_inp <= "000000000000000000011000011101100101" else
--"0000010111111101" when sig_inp <= "000000000000000000011000011111110110" else
--"0000010111110110" when sig_inp <= "000000000000000000011000100010001000" else
--"0000010111101111" when sig_inp <= "000000000000000000011000100100011010" else
--"0000010111101000" when sig_inp <= "000000000000000000011000100110101011" else
--"0000010111100001" when sig_inp <= "000000000000000000011000101000111101" else
--"0000010111011011" when sig_inp <= "000000000000000000011000101011001111" else
--"0000010111010100" when sig_inp <= "000000000000000000011000101101100000" else
--"0000010111001110" when sig_inp <= "000000000000000000011000101111110010" else
--"0000010111000111" when sig_inp <= "000000000000000000011000110010000011" else
--"0000010111000000" when sig_inp <= "000000000000000000011000110100010101" else
--"0000010110111010" when sig_inp <= "000000000000000000011000110110100111" else
--"0000010110110011" when sig_inp <= "000000000000000000011000111000111000" else
--"0000010110101101" when sig_inp <= "000000000000000000011000111011001010" else
--"0000010110100110" when sig_inp <= "000000000000000000011000111101011100" else
--"0000010110100000" when sig_inp <= "000000000000000000011000111111101101" else
--"0000010110011010" when sig_inp <= "000000000000000000011001000001111111" else
--"0000010110010011" when sig_inp <= "000000000000000000011001000100010001" else
--"0000010110001101" when sig_inp <= "000000000000000000011001000110100010" else
--"0000010110000111" when sig_inp <= "000000000000000000011001001000110100" else
--"0000010110000000" when sig_inp <= "000000000000000000011001001011000101" else
--"0000010101111010" when sig_inp <= "000000000000000000011001001101010111" else
--"0000010101110100" when sig_inp <= "000000000000000000011001001111101001" else
--"0000010101101110" when sig_inp <= "000000000000000000011001010001111010" else
--"0000010101101000" when sig_inp <= "000000000000000000011001010100001100" else
--"0000010101100001" when sig_inp <= "000000000000000000011001010110011110" else
--"0000010101011011" when sig_inp <= "000000000000000000011001011000101111" else
--"0000010101010101" when sig_inp <= "000000000000000000011001011011000001" else
--"0000010101001111" when sig_inp <= "000000000000000000011001011101010011" else
--"0000010101001001" when sig_inp <= "000000000000000000011001011111100100" else
--"0000010101000011" when sig_inp <= "000000000000000000011001100001110110" else
--"0000010100111101" when sig_inp <= "000000000000000000011001100100000111" else
--"0000010100110111" when sig_inp <= "000000000000000000011001100110011001" else
--"0000010100110001" when sig_inp <= "000000000000000000011001101000101011" else
--"0000010100101011" when sig_inp <= "000000000000000000011001101010111100" else
--"0000010100100110" when sig_inp <= "000000000000000000011001101101001110" else
--"0000010100100000" when sig_inp <= "000000000000000000011001101111100000" else
--"0000010100011010" when sig_inp <= "000000000000000000011001110001110001" else
--"0000010100010100" when sig_inp <= "000000000000000000011001110100000011" else
--"0000010100001110" when sig_inp <= "000000000000000000011001110110010101" else
--"0000010100001001" when sig_inp <= "000000000000000000011001111000100110" else
--"0000010100000011" when sig_inp <= "000000000000000000011001111010111000" else
--"0000010011111101" when sig_inp <= "000000000000000000011001111101001001" else
--"0000010011110111" when sig_inp <= "000000000000000000011001111111011011" else
--"0000010011110010" when sig_inp <= "000000000000000000011010000001101101" else
--"0000010011101100" when sig_inp <= "000000000000000000011010000011111110" else
--"0000010011100111" when sig_inp <= "000000000000000000011010000110010000" else
--"0000010011100001" when sig_inp <= "000000000000000000011010001000100010" else
--"0000010011011100" when sig_inp <= "000000000000000000011010001010110011" else
--"0000010011010110" when sig_inp <= "000000000000000000011010001101000101" else
--"0000010011010001" when sig_inp <= "000000000000000000011010001111010111" else
--"0000010011001011" when sig_inp <= "000000000000000000011010010001101000" else
--"0000010011000110" when sig_inp <= "000000000000000000011010010011111010" else
--"0000010011000000" when sig_inp <= "000000000000000000011010010110001011" else
--"0000010010111011" when sig_inp <= "000000000000000000011010011000011101" else
--"0000010010110101" when sig_inp <= "000000000000000000011010011010101111" else
--"0000010010110000" when sig_inp <= "000000000000000000011010011101000000" else
--"0000010010101011" when sig_inp <= "000000000000000000011010011111010010" else
--"0000010010100101" when sig_inp <= "000000000000000000011010100001100100" else
--"0000010010100000" when sig_inp <= "000000000000000000011010100011110101" else
--"0000010010011011" when sig_inp <= "000000000000000000011010100110000111" else
--"0000010010010110" when sig_inp <= "000000000000000000011010101000011001" else
--"0000010010010000" when sig_inp <= "000000000000000000011010101010101010" else
--"0000010010001011" when sig_inp <= "000000000000000000011010101100111100" else
--"0000010010000110" when sig_inp <= "000000000000000000011010101111001101" else
--"0000010010000001" when sig_inp <= "000000000000000000011010110001011111" else
--"0000010001111100" when sig_inp <= "000000000000000000011010110011110001" else
--"0000010001110111" when sig_inp <= "000000000000000000011010110110000010" else
--"0000010001110010" when sig_inp <= "000000000000000000011010111000010100" else
--"0000010001101101" when sig_inp <= "000000000000000000011010111010100110" else
--"0000010001101000" when sig_inp <= "000000000000000000011010111100110111" else
--"0000010001100011" when sig_inp <= "000000000000000000011010111111001001" else
--"0000010001011110" when sig_inp <= "000000000000000000011011000001011011" else
--"0000010001011001" when sig_inp <= "000000000000000000011011000011101100" else
--"0000010001010100" when sig_inp <= "000000000000000000011011000101111110" else
--"0000010001001111" when sig_inp <= "000000000000000000011011001000001111" else
--"0000010001001010" when sig_inp <= "000000000000000000011011001010100001" else
--"0000010001000101" when sig_inp <= "000000000000000000011011001100110011" else
--"0000010001000000" when sig_inp <= "000000000000000000011011001111000100" else
--"0000010000111011" when sig_inp <= "000000000000000000011011010001010110" else
--"0000010000110111" when sig_inp <= "000000000000000000011011010011101000" else
--"0000010000110010" when sig_inp <= "000000000000000000011011010101111001" else
--"0000010000101101" when sig_inp <= "000000000000000000011011011000001011" else
--"0000010000101000" when sig_inp <= "000000000000000000011011011010011101" else
--"0000010000100100" when sig_inp <= "000000000000000000011011011100101110" else
--"0000010000011111" when sig_inp <= "000000000000000000011011011111000000" else
--"0000010000011010" when sig_inp <= "000000000000000000011011100001010001" else
--"0000010000010110" when sig_inp <= "000000000000000000011011100011100011" else
--"0000010000010001" when sig_inp <= "000000000000000000011011100101110101" else
--"0000010000001100" when sig_inp <= "000000000000000000011011101000000110" else
--"0000010000001000" when sig_inp <= "000000000000000000011011101010011000" else
--"0000010000000011" when sig_inp <= "000000000000000000011011101100101010" else
--"0000001111111111" when sig_inp <= "000000000000000000011011101110111011" else
--"0000001111111010" when sig_inp <= "000000000000000000011011110001001101" else
--"0000001111110101" when sig_inp <= "000000000000000000011011110011011111" else
--"0000001111110001" when sig_inp <= "000000000000000000011011110101110000" else
--"0000001111101101" when sig_inp <= "000000000000000000011011111000000010" else
--"0000001111101000" when sig_inp <= "000000000000000000011011111010010011" else
--"0000001111100100" when sig_inp <= "000000000000000000011011111100100101" else
--"0000001111011111" when sig_inp <= "000000000000000000011011111110110111" else
--"0000001111011011" when sig_inp <= "000000000000000000011100000001001000" else
--"0000001111010110" when sig_inp <= "000000000000000000011100000011011010" else
--"0000001111010010" when sig_inp <= "000000000000000000011100000101101100" else
--"0000001111001110" when sig_inp <= "000000000000000000011100000111111101" else
--"0000001111001001" when sig_inp <= "000000000000000000011100001010001111" else
--"0000001111000101" when sig_inp <= "000000000000000000011100001100100000" else
--"0000001111000001" when sig_inp <= "000000000000000000011100001110110010" else
--"0000001110111101" when sig_inp <= "000000000000000000011100010001000100" else
--"0000001110111000" when sig_inp <= "000000000000000000011100010011010101" else
--"0000001110110100" when sig_inp <= "000000000000000000011100010101100111" else
--"0000001110110000" when sig_inp <= "000000000000000000011100010111111001" else
--"0000001110101100" when sig_inp <= "000000000000000000011100011010001010" else
--"0000001110101000" when sig_inp <= "000000000000000000011100011100011100" else
--"0000001110100011" when sig_inp <= "000000000000000000011100011110101110" else
--"0000001110011111" when sig_inp <= "000000000000000000011100100000111111" else
--"0000001110011011" when sig_inp <= "000000000000000000011100100011010001" else
--"0000001110010111" when sig_inp <= "000000000000000000011100100101100010" else
--"0000001110010011" when sig_inp <= "000000000000000000011100100111110100" else
--"0000001110001111" when sig_inp <= "000000000000000000011100101010000110" else
--"0000001110001011" when sig_inp <= "000000000000000000011100101100010111" else
--"0000001110000111" when sig_inp <= "000000000000000000011100101110101001" else
--"0000001110000011" when sig_inp <= "000000000000000000011100110000111011" else
--"0000001101111111" when sig_inp <= "000000000000000000011100110011001100" else
--"0000001101111011" when sig_inp <= "000000000000000000011100110101011110" else
--"0000001101110111" when sig_inp <= "000000000000000000011100110111110000" else
--"0000001101110011" when sig_inp <= "000000000000000000011100111010000001" else
--"0000001101101111" when sig_inp <= "000000000000000000011100111100010011" else
--"0000001101101011" when sig_inp <= "000000000000000000011100111110100100" else
--"0000001101100111" when sig_inp <= "000000000000000000011101000000110110" else
--"0000001101100011" when sig_inp <= "000000000000000000011101000011001000" else
--"0000001101100000" when sig_inp <= "000000000000000000011101000101011001" else
--"0000001101011100" when sig_inp <= "000000000000000000011101000111101011" else
--"0000001101011000" when sig_inp <= "000000000000000000011101001001111101" else
--"0000001101010100" when sig_inp <= "000000000000000000011101001100001110" else
--"0000001101010000" when sig_inp <= "000000000000000000011101001110100000" else
--"0000001101001101" when sig_inp <= "000000000000000000011101010000110010" else
--"0000001101001001" when sig_inp <= "000000000000000000011101010011000011" else
--"0000001101000101" when sig_inp <= "000000000000000000011101010101010101" else
--"0000001101000001" when sig_inp <= "000000000000000000011101010111100110" else
--"0000001100111110" when sig_inp <= "000000000000000000011101011001111000" else
--"0000001100111010" when sig_inp <= "000000000000000000011101011100001010" else
--"0000001100110110" when sig_inp <= "000000000000000000011101011110011011" else
--"0000001100110011" when sig_inp <= "000000000000000000011101100000101101" else
--"0000001100101111" when sig_inp <= "000000000000000000011101100010111111" else
--"0000001100101011" when sig_inp <= "000000000000000000011101100101010000" else
--"0000001100101000" when sig_inp <= "000000000000000000011101100111100010" else
--"0000001100100100" when sig_inp <= "000000000000000000011101101001110100" else
--"0000001100100001" when sig_inp <= "000000000000000000011101101100000101" else
--"0000001100011101" when sig_inp <= "000000000000000000011101101110010111" else
--"0000001100011010" when sig_inp <= "000000000000000000011101110000101000" else
--"0000001100010110" when sig_inp <= "000000000000000000011101110010111010" else
--"0000001100010011" when sig_inp <= "000000000000000000011101110101001100" else
--"0000001100001111" when sig_inp <= "000000000000000000011101110111011101" else
--"0000001100001100" when sig_inp <= "000000000000000000011101111001101111" else
--"0000001100001000" when sig_inp <= "000000000000000000011101111100000001" else
--"0000001100000101" when sig_inp <= "000000000000000000011101111110010010" else
--"0000001100000001" when sig_inp <= "000000000000000000011110000000100100" else
--"0000001011111110" when sig_inp <= "000000000000000000011110000010110110" else
--"0000001011111010" when sig_inp <= "000000000000000000011110000101000111" else
--"0000001011110111" when sig_inp <= "000000000000000000011110000111011001" else
--"0000001011110100" when sig_inp <= "000000000000000000011110001001101010" else
--"0000001011110000" when sig_inp <= "000000000000000000011110001011111100" else
--"0000001011101101" when sig_inp <= "000000000000000000011110001110001110" else
--"0000001011101010" when sig_inp <= "000000000000000000011110010000011111" else
--"0000001011100110" when sig_inp <= "000000000000000000011110010010110001" else
--"0000001011100011" when sig_inp <= "000000000000000000011110010101000011" else
--"0000001011100000" when sig_inp <= "000000000000000000011110010111010100" else
--"0000001011011101" when sig_inp <= "000000000000000000011110011001100110" else
--"0000001011011001" when sig_inp <= "000000000000000000011110011011111000" else
--"0000001011010110" when sig_inp <= "000000000000000000011110011110001001" else
--"0000001011010011" when sig_inp <= "000000000000000000011110100000011011" else
--"0000001011010000" when sig_inp <= "000000000000000000011110100010101100" else
--"0000001011001100" when sig_inp <= "000000000000000000011110100100111110" else
--"0000001011001001" when sig_inp <= "000000000000000000011110100111010000" else
--"0000001011000110" when sig_inp <= "000000000000000000011110101001100001" else
--"0000001011000011" when sig_inp <= "000000000000000000011110101011110011" else
--"0000001011000000" when sig_inp <= "000000000000000000011110101110000101" else
--"0000001010111101" when sig_inp <= "000000000000000000011110110000010110" else
--"0000001010111010" when sig_inp <= "000000000000000000011110110010101000" else
--"0000001010110110" when sig_inp <= "000000000000000000011110110100111010" else
--"0000001010110011" when sig_inp <= "000000000000000000011110110111001011" else
--"0000001010110000" when sig_inp <= "000000000000000000011110111001011101" else
--"0000001010101101" when sig_inp <= "000000000000000000011110111011101110" else
--"0000001010101010" when sig_inp <= "000000000000000000011110111110000000" else
--"0000001010100111" when sig_inp <= "000000000000000000011111000000010010" else
--"0000001010100100" when sig_inp <= "000000000000000000011111000010100011" else
--"0000001010100001" when sig_inp <= "000000000000000000011111000100110101" else
--"0000001010011110" when sig_inp <= "000000000000000000011111000111000111" else
--"0000001010011011" when sig_inp <= "000000000000000000011111001001011000" else
--"0000001010011000" when sig_inp <= "000000000000000000011111001011101010" else
--"0000001010010101" when sig_inp <= "000000000000000000011111001101111100" else
--"0000001010010010" when sig_inp <= "000000000000000000011111010000001101" else
--"0000001010001111" when sig_inp <= "000000000000000000011111010010011111" else
--"0000001010001101" when sig_inp <= "000000000000000000011111010100110000" else
--"0000001010001010" when sig_inp <= "000000000000000000011111010111000010" else
--"0000001010000111" when sig_inp <= "000000000000000000011111011001010100" else
--"0000001010000100" when sig_inp <= "000000000000000000011111011011100101" else
--"0000001010000001" when sig_inp <= "000000000000000000011111011101110111" else
--"0000001001111110" when sig_inp <= "000000000000000000011111100000001001" else
--"0000001001111011" when sig_inp <= "000000000000000000011111100010011010" else
--"0000001001111001" when sig_inp <= "000000000000000000011111100100101100" else
--"0000001001110110" when sig_inp <= "000000000000000000011111100110111110" else
--"0000001001110011" when sig_inp <= "000000000000000000011111101001001111" else
--"0000001001110000" when sig_inp <= "000000000000000000011111101011100001" else
--"0000001001101101" when sig_inp <= "000000000000000000011111101101110010" else
--"0000001001101011" when sig_inp <= "000000000000000000011111110000000100" else
--"0000001001101000" when sig_inp <= "000000000000000000011111110010010110" else
--"0000001001100101" when sig_inp <= "000000000000000000011111110100100111" else
--"0000001001100010" when sig_inp <= "000000000000000000011111110110111001" else
--"0000001001100000" when sig_inp <= "000000000000000000011111111001001011" else
--"0000001001011101" when sig_inp <= "000000000000000000011111111011011100" else
--"0000001001011010" when sig_inp <= "000000000000000000011111111101101110" else
--"0000001001011000" when sig_inp <= "000000000000000000100000000000000000" else
--"0000001001010101" when sig_inp <= "000000000000000000100000000010010001" else
--"0000001001010010" when sig_inp <= "000000000000000000100000000100100011" else
--"0000001001010000" when sig_inp <= "000000000000000000100000000110110100" else
--"0000001001001101" when sig_inp <= "000000000000000000100000001001000110" else
--"0000001001001010" when sig_inp <= "000000000000000000100000001011011000" else
--"0000001001001000" when sig_inp <= "000000000000000000100000001101101001" else
--"0000001001000101" when sig_inp <= "000000000000000000100000001111111011" else
--"0000001001000011" when sig_inp <= "000000000000000000100000010010001101" else
--"0000001001000000" when sig_inp <= "000000000000000000100000010100011110" else
--"0000001000111110" when sig_inp <= "000000000000000000100000010110110000" else
--"0000001000111011" when sig_inp <= "000000000000000000100000011001000001" else
--"0000001000111000" when sig_inp <= "000000000000000000100000011011010011" else
--"0000001000110110" when sig_inp <= "000000000000000000100000011101100101" else
--"0000001000110011" when sig_inp <= "000000000000000000100000011111110110" else
--"0000001000110001" when sig_inp <= "000000000000000000100000100010001000" else
--"0000001000101110" when sig_inp <= "000000000000000000100000100100011010" else
--"0000001000101100" when sig_inp <= "000000000000000000100000100110101011" else
--"0000001000101010" when sig_inp <= "000000000000000000100000101000111101" else
--"0000001000100111" when sig_inp <= "000000000000000000100000101011001111" else
--"0000001000100101" when sig_inp <= "000000000000000000100000101101100000" else
--"0000001000100010" when sig_inp <= "000000000000000000100000101111110010" else
--"0000001000100000" when sig_inp <= "000000000000000000100000110010000011" else
--"0000001000011101" when sig_inp <= "000000000000000000100000110100010101" else
--"0000001000011011" when sig_inp <= "000000000000000000100000110110100111" else
--"0000001000011001" when sig_inp <= "000000000000000000100000111000111000" else
--"0000001000010110" when sig_inp <= "000000000000000000100000111011001010" else
--"0000001000010100" when sig_inp <= "000000000000000000100000111101011100" else
--"0000001000010001" when sig_inp <= "000000000000000000100000111111101101" else
--"0000001000001111" when sig_inp <= "000000000000000000100001000001111111" else
--"0000001000001101" when sig_inp <= "000000000000000000100001000100010001" else
--"0000001000001010" when sig_inp <= "000000000000000000100001000110100010" else
--"0000001000001000" when sig_inp <= "000000000000000000100001001000110100" else
--"0000001000000110" when sig_inp <= "000000000000000000100001001011000101" else
--"0000001000000011" when sig_inp <= "000000000000000000100001001101010111" else
--"0000001000000001" when sig_inp <= "000000000000000000100001001111101001" else
--"0000000111111111" when sig_inp <= "000000000000000000100001010001111010" else
--"0000000111111101" when sig_inp <= "000000000000000000100001010100001100" else
--"0000000111111010" when sig_inp <= "000000000000000000100001010110011110" else
--"0000000111111000" when sig_inp <= "000000000000000000100001011000101111" else
--"0000000111110110" when sig_inp <= "000000000000000000100001011011000001" else
--"0000000111110100" when sig_inp <= "000000000000000000100001011101010011" else
--"0000000111110001" when sig_inp <= "000000000000000000100001011111100100" else
--"0000000111101111" when sig_inp <= "000000000000000000100001100001110110" else
--"0000000111101101" when sig_inp <= "000000000000000000100001100100000111" else
--"0000000111101011" when sig_inp <= "000000000000000000100001100110011001" else
--"0000000111101001" when sig_inp <= "000000000000000000100001101000101011" else
--"0000000111100111" when sig_inp <= "000000000000000000100001101010111100" else
--"0000000111100100" when sig_inp <= "000000000000000000100001101101001110" else
--"0000000111100010" when sig_inp <= "000000000000000000100001101111100000" else
--"0000000111100000" when sig_inp <= "000000000000000000100001110001110001" else
--"0000000111011110" when sig_inp <= "000000000000000000100001110100000011" else
--"0000000111011100" when sig_inp <= "000000000000000000100001110110010101" else
--"0000000111011010" when sig_inp <= "000000000000000000100001111000100110" else
--"0000000111011000" when sig_inp <= "000000000000000000100001111010111000" else
--"0000000111010110" when sig_inp <= "000000000000000000100001111101001001" else
--"0000000111010011" when sig_inp <= "000000000000000000100001111111011011" else
--"0000000111010001" when sig_inp <= "000000000000000000100010000001101101" else
--"0000000111001111" when sig_inp <= "000000000000000000100010000011111110" else
--"0000000111001101" when sig_inp <= "000000000000000000100010000110010000" else
--"0000000111001011" when sig_inp <= "000000000000000000100010001000100010" else
--"0000000111001001" when sig_inp <= "000000000000000000100010001010110011" else
--"0000000111000111" when sig_inp <= "000000000000000000100010001101000101" else
--"0000000111000101" when sig_inp <= "000000000000000000100010001111010111" else
--"0000000111000011" when sig_inp <= "000000000000000000100010010001101000" else
--"0000000111000001" when sig_inp <= "000000000000000000100010010011111010" else
--"0000000110111111" when sig_inp <= "000000000000000000100010010110001011" else
--"0000000110111101" when sig_inp <= "000000000000000000100010011000011101" else
--"0000000110111011" when sig_inp <= "000000000000000000100010011010101111" else
--"0000000110111001" when sig_inp <= "000000000000000000100010011101000000" else
--"0000000110110111" when sig_inp <= "000000000000000000100010011111010010" else
--"0000000110110101" when sig_inp <= "000000000000000000100010100001100100" else
--"0000000110110011" when sig_inp <= "000000000000000000100010100011110101" else
--"0000000110110001" when sig_inp <= "000000000000000000100010100110000111" else
--"0000000110101111" when sig_inp <= "000000000000000000100010101000011001" else
--"0000000110101110" when sig_inp <= "000000000000000000100010101010101010" else
--"0000000110101100" when sig_inp <= "000000000000000000100010101100111100" else
--"0000000110101010" when sig_inp <= "000000000000000000100010101111001101" else
--"0000000110101000" when sig_inp <= "000000000000000000100010110001011111" else
--"0000000110100110" when sig_inp <= "000000000000000000100010110011110001" else
--"0000000110100100" when sig_inp <= "000000000000000000100010110110000010" else
--"0000000110100010" when sig_inp <= "000000000000000000100010111000010100" else
--"0000000110100000" when sig_inp <= "000000000000000000100010111010100110" else
--"0000000110011111" when sig_inp <= "000000000000000000100010111100110111" else
--"0000000110011101" when sig_inp <= "000000000000000000100010111111001001" else
--"0000000110011011" when sig_inp <= "000000000000000000100011000001011011" else
--"0000000110011001" when sig_inp <= "000000000000000000100011000011101100" else
--"0000000110010111" when sig_inp <= "000000000000000000100011000101111110" else
--"0000000110010101" when sig_inp <= "000000000000000000100011001000001111" else
--"0000000110010100" when sig_inp <= "000000000000000000100011001010100001" else
--"0000000110010010" when sig_inp <= "000000000000000000100011001100110011" else
--"0000000110010000" when sig_inp <= "000000000000000000100011001111000100" else
--"0000000110001110" when sig_inp <= "000000000000000000100011010001010110" else
--"0000000110001100" when sig_inp <= "000000000000000000100011010011101000" else
--"0000000110001011" when sig_inp <= "000000000000000000100011010101111001" else
--"0000000110001001" when sig_inp <= "000000000000000000100011011000001011" else
--"0000000110000111" when sig_inp <= "000000000000000000100011011010011101" else
--"0000000110000101" when sig_inp <= "000000000000000000100011011100101110" else
--"0000000110000100" when sig_inp <= "000000000000000000100011011111000000" else
--"0000000110000010" when sig_inp <= "000000000000000000100011100001010001" else
--"0000000110000000" when sig_inp <= "000000000000000000100011100011100011" else
--"0000000101111111" when sig_inp <= "000000000000000000100011100101110101" else
--"0000000101111101" when sig_inp <= "000000000000000000100011101000000110" else
--"0000000101111011" when sig_inp <= "000000000000000000100011101010011000" else
--"0000000101111010" when sig_inp <= "000000000000000000100011101100101010" else
--"0000000101111000" when sig_inp <= "000000000000000000100011101110111011" else
--"0000000101110110" when sig_inp <= "000000000000000000100011110001001101" else
--"0000000101110101" when sig_inp <= "000000000000000000100011110011011111" else
--"0000000101110011" when sig_inp <= "000000000000000000100011110101110000" else
--"0000000101110001" when sig_inp <= "000000000000000000100011111000000010" else
--"0000000101110000" when sig_inp <= "000000000000000000100011111010010011" else
--"0000000101101110" when sig_inp <= "000000000000000000100011111100100101" else
--"0000000101101100" when sig_inp <= "000000000000000000100011111110110111" else
--"0000000101101011" when sig_inp <= "000000000000000000100100000001001000" else
--"0000000101101001" when sig_inp <= "000000000000000000100100000011011010" else
--"0000000101100111" when sig_inp <= "000000000000000000100100000101101100" else
--"0000000101100110" when sig_inp <= "000000000000000000100100000111111101" else
--"0000000101100100" when sig_inp <= "000000000000000000100100001010001111" else
--"0000000101100011" when sig_inp <= "000000000000000000100100001100100000" else
--"0000000101100001" when sig_inp <= "000000000000000000100100001110110010" else
--"0000000101100000" when sig_inp <= "000000000000000000100100010001000100" else
--"0000000101011110" when sig_inp <= "000000000000000000100100010011010101" else
--"0000000101011100" when sig_inp <= "000000000000000000100100010101100111" else
--"0000000101011011" when sig_inp <= "000000000000000000100100010111111001" else
--"0000000101011001" when sig_inp <= "000000000000000000100100011010001010" else
--"0000000101011000" when sig_inp <= "000000000000000000100100011100011100" else
--"0000000101010110" when sig_inp <= "000000000000000000100100011110101110" else
--"0000000101010101" when sig_inp <= "000000000000000000100100100000111111" else
--"0000000101010011" when sig_inp <= "000000000000000000100100100011010001" else
--"0000000101010010" when sig_inp <= "000000000000000000100100100101100010" else
--"0000000101010000" when sig_inp <= "000000000000000000100100100111110100" else
--"0000000101001111" when sig_inp <= "000000000000000000100100101010000110" else
--"0000000101001101" when sig_inp <= "000000000000000000100100101100010111" else
--"0000000101001100" when sig_inp <= "000000000000000000100100101110101001" else
--"0000000101001010" when sig_inp <= "000000000000000000100100110000111011" else
--"0000000101001001" when sig_inp <= "000000000000000000100100110011001100" else
--"0000000101000111" when sig_inp <= "000000000000000000100100110101011110" else
--"0000000101000110" when sig_inp <= "000000000000000000100100110111110000" else
--"0000000101000101" when sig_inp <= "000000000000000000100100111010000001" else
--"0000000101000011" when sig_inp <= "000000000000000000100100111100010011" else
--"0000000101000010" when sig_inp <= "000000000000000000100100111110100100" else
--"0000000101000000" when sig_inp <= "000000000000000000100101000000110110" else
--"0000000100111111" when sig_inp <= "000000000000000000100101000011001000" else
--"0000000100111101" when sig_inp <= "000000000000000000100101000101011001" else
--"0000000100111100" when sig_inp <= "000000000000000000100101000111101011" else
--"0000000100111011" when sig_inp <= "000000000000000000100101001001111101" else
--"0000000100111001" when sig_inp <= "000000000000000000100101001100001110" else
--"0000000100111000" when sig_inp <= "000000000000000000100101001110100000" else
--"0000000100110110" when sig_inp <= "000000000000000000100101010000110010" else
--"0000000100110101" when sig_inp <= "000000000000000000100101010011000011" else
--"0000000100110100" when sig_inp <= "000000000000000000100101010101010101" else
--"0000000100110010" when sig_inp <= "000000000000000000100101010111100110" else
--"0000000100110001" when sig_inp <= "000000000000000000100101011001111000" else
--"0000000100110000" when sig_inp <= "000000000000000000100101011100001010" else
--"0000000100101110" when sig_inp <= "000000000000000000100101011110011011" else
--"0000000100101101" when sig_inp <= "000000000000000000100101100000101101" else
--"0000000100101100" when sig_inp <= "000000000000000000100101100010111111" else
--"0000000100101010" when sig_inp <= "000000000000000000100101100101010000" else
--"0000000100101001" when sig_inp <= "000000000000000000100101100111100010" else
--"0000000100101000" when sig_inp <= "000000000000000000100101101001110100" else
--"0000000100100110" when sig_inp <= "000000000000000000100101101100000101" else
--"0000000100100101" when sig_inp <= "000000000000000000100101101110010111" else
--"0000000100100100" when sig_inp <= "000000000000000000100101110000101000" else
--"0000000100100010" when sig_inp <= "000000000000000000100101110010111010" else
--"0000000100100001" when sig_inp <= "000000000000000000100101110101001100" else
--"0000000100100000" when sig_inp <= "000000000000000000100101110111011101" else
--"0000000100011110" when sig_inp <= "000000000000000000100101111001101111" else
--"0000000100011101" when sig_inp <= "000000000000000000100101111100000001" else
--"0000000100011100" when sig_inp <= "000000000000000000100101111110010010" else
--"0000000100011011" when sig_inp <= "000000000000000000100110000000100100" else
--"0000000100011001" when sig_inp <= "000000000000000000100110000010110110" else
--"0000000100011000" when sig_inp <= "000000000000000000100110000101000111" else
--"0000000100010111" when sig_inp <= "000000000000000000100110000111011001" else
--"0000000100010110" when sig_inp <= "000000000000000000100110001001101010" else
--"0000000100010100" when sig_inp <= "000000000000000000100110001011111100" else
--"0000000100010011" when sig_inp <= "000000000000000000100110001110001110" else
--"0000000100010010" when sig_inp <= "000000000000000000100110010000011111" else
--"0000000100010001" when sig_inp <= "000000000000000000100110010010110001" else
--"0000000100010000" when sig_inp <= "000000000000000000100110010101000011" else
--"0000000100001110" when sig_inp <= "000000000000000000100110010111010100" else
--"0000000100001101" when sig_inp <= "000000000000000000100110011001100110" else
--"0000000100001100" when sig_inp <= "000000000000000000100110011011111000" else
--"0000000100001011" when sig_inp <= "000000000000000000100110011110001001" else
--"0000000100001010" when sig_inp <= "000000000000000000100110100000011011" else
--"0000000100001000" when sig_inp <= "000000000000000000100110100010101100" else
--"0000000100000111" when sig_inp <= "000000000000000000100110100100111110" else
--"0000000100000110" when sig_inp <= "000000000000000000100110100111010000" else
--"0000000100000101" when sig_inp <= "000000000000000000100110101001100001" else
--"0000000100000100" when sig_inp <= "000000000000000000100110101011110011" else
--"0000000100000011" when sig_inp <= "000000000000000000100110101110000101" else
--"0000000100000001" when sig_inp <= "000000000000000000100110110000010110" else
--"0000000100000000" when sig_inp <= "000000000000000000100110110010101000" else
--"0000000011111111" when sig_inp <= "000000000000000000100110110100111010" else
--"0000000011111110" when sig_inp <= "000000000000000000100110110111001011" else
--"0000000011111101" when sig_inp <= "000000000000000000100110111001011101" else
--"0000000011111100" when sig_inp <= "000000000000000000100110111011101110" else
--"0000000011111011" when sig_inp <= "000000000000000000100110111110000000" else
--"0000000011111010" when sig_inp <= "000000000000000000100111000000010010" else
--"0000000011111000" when sig_inp <= "000000000000000000100111000010100011" else
--"0000000011110111" when sig_inp <= "000000000000000000100111000100110101" else
--"0000000011110110" when sig_inp <= "000000000000000000100111000111000111" else
--"0000000011110101" when sig_inp <= "000000000000000000100111001001011000" else
--"0000000011110100" when sig_inp <= "000000000000000000100111001011101010" else
--"0000000011110011" when sig_inp <= "000000000000000000100111001101111100" else
--"0000000011110010" when sig_inp <= "000000000000000000100111010000001101" else
--"0000000011110001" when sig_inp <= "000000000000000000100111010010011111" else
--"0000000011110000" when sig_inp <= "000000000000000000100111010100110000" else
--"0000000011101111" when sig_inp <= "000000000000000000100111010111000010" else
--"0000000011101110" when sig_inp <= "000000000000000000100111011001010100" else
--"0000000011101101" when sig_inp <= "000000000000000000100111011011100101" else
--"0000000011101100" when sig_inp <= "000000000000000000100111011101110111" else
--"0000000011101010" when sig_inp <= "000000000000000000100111100000001001" else
--"0000000011101001" when sig_inp <= "000000000000000000100111100010011010" else
--"0000000011101000" when sig_inp <= "000000000000000000100111100100101100" else
--"0000000011100111" when sig_inp <= "000000000000000000100111100110111110" else
--"0000000011100110" when sig_inp <= "000000000000000000100111101001001111" else
--"0000000011100101" when sig_inp <= "000000000000000000100111101011100001" else
--"0000000011100100" when sig_inp <= "000000000000000000100111101101110010" else
--"0000000011100011" when sig_inp <= "000000000000000000100111110000000100" else
--"0000000011100010" when sig_inp <= "000000000000000000100111110010010110" else
--"0000000011100001" when sig_inp <= "000000000000000000100111110100100111" else
--"0000000011100000" when sig_inp <= "000000000000000000100111110110111001" else
--"0000000011011111" when sig_inp <= "000000000000000000100111111001001011" else
--"0000000011011110" when sig_inp <= "000000000000000000100111111011011100" else
--"0000000011011101" when sig_inp <= "000000000000000000100111111101101110" else
--"0000000011011100" when sig_inp <= "000000000000000000101000000000000000" else
--"0000000011011011" when sig_inp <= "000000000000000000101000000010010001" else
--"0000000011011010" when sig_inp <= "000000000000000000101000000100100011" else
--"0000000011011001" when sig_inp <= "000000000000000000101000000110110100" else
--"0000000011011000" when sig_inp <= "000000000000000000101000001001000110" else
--"0000000011010111" when sig_inp <= "000000000000000000101000001011011000" else
--"0000000011010110" when sig_inp <= "000000000000000000101000001101101001" else
--"0000000011010101" when sig_inp <= "000000000000000000101000010010001101" else
--"0000000011010100" when sig_inp <= "000000000000000000101000010100011110" else
--"0000000011010011" when sig_inp <= "000000000000000000101000010110110000" else
--"0000000011010010" when sig_inp <= "000000000000000000101000011001000001" else
--"0000000011010001" when sig_inp <= "000000000000000000101000011011010011" else
--"0000000011010000" when sig_inp <= "000000000000000000101000011101100101" else
--"0000000011001111" when sig_inp <= "000000000000000000101000011111110110" else
--"0000000011001110" when sig_inp <= "000000000000000000101000100010001000" else
--"0000000011001101" when sig_inp <= "000000000000000000101000100100011010" else
--"0000000011001100" when sig_inp <= "000000000000000000101000100110101011" else
--"0000000011001011" when sig_inp <= "000000000000000000101000101000111101" else
--"0000000011001010" when sig_inp <= "000000000000000000101000101011001111" else
--"0000000011001001" when sig_inp <= "000000000000000000101000101111110010" else
--"0000000011001000" when sig_inp <= "000000000000000000101000110010000011" else
--"0000000011000111" when sig_inp <= "000000000000000000101000110100010101" else
--"0000000011000110" when sig_inp <= "000000000000000000101000110110100111" else
--"0000000011000101" when sig_inp <= "000000000000000000101000111000111000" else
--"0000000011000100" when sig_inp <= "000000000000000000101000111011001010" else
--"0000000011000011" when sig_inp <= "000000000000000000101000111101011100" else
--"0000000011000010" when sig_inp <= "000000000000000000101000111111101101" else
--"0000000011000001" when sig_inp <= "000000000000000000101001000100010001" else
--"0000000011000000" when sig_inp <= "000000000000000000101001000110100010" else
--"0000000010111111" when sig_inp <= "000000000000000000101001001000110100" else
--"0000000010111110" when sig_inp <= "000000000000000000101001001011000101" else
--"0000000010111101" when sig_inp <= "000000000000000000101001001101010111" else
--"0000000010111100" when sig_inp <= "000000000000000000101001001111101001" else
--"0000000010111011" when sig_inp <= "000000000000000000101001010100001100" else
--"0000000010111010" when sig_inp <= "000000000000000000101001010110011110" else
--"0000000010111001" when sig_inp <= "000000000000000000101001011000101111" else
--"0000000010111000" when sig_inp <= "000000000000000000101001011011000001" else
--"0000000010110111" when sig_inp <= "000000000000000000101001011111100100" else
--"0000000010110110" when sig_inp <= "000000000000000000101001100001110110" else
--"0000000010110101" when sig_inp <= "000000000000000000101001100100000111" else
--"0000000010110100" when sig_inp <= "000000000000000000101001100110011001" else
--"0000000010110011" when sig_inp <= "000000000000000000101001101000101011" else
--"0000000010110010" when sig_inp <= "000000000000000000101001101101001110" else
--"0000000010110001" when sig_inp <= "000000000000000000101001101111100000" else
--"0000000010110000" when sig_inp <= "000000000000000000101001110001110001" else
--"0000000010101111" when sig_inp <= "000000000000000000101001110110010101" else
--"0000000010101110" when sig_inp <= "000000000000000000101001111000100110" else
--"0000000010101101" when sig_inp <= "000000000000000000101001111010111000" else
--"0000000010101100" when sig_inp <= "000000000000000000101001111101001001" else
--"0000000010101011" when sig_inp <= "000000000000000000101010000001101101" else
--"0000000010101010" when sig_inp <= "000000000000000000101010000011111110" else
--"0000000010101001" when sig_inp <= "000000000000000000101010000110010000" else
--"0000000010101000" when sig_inp <= "000000000000000000101010001010110011" else
--"0000000010100111" when sig_inp <= "000000000000000000101010001101000101" else
--"0000000010100110" when sig_inp <= "000000000000000000101010001111010111" else
--"0000000010100101" when sig_inp <= "000000000000000000101010010011111010" else
--"0000000010100100" when sig_inp <= "000000000000000000101010010110001011" else
--"0000000010100011" when sig_inp <= "000000000000000000101010011000011101" else
--"0000000010100010" when sig_inp <= "000000000000000000101010011101000000" else
--"0000000010100001" when sig_inp <= "000000000000000000101010011111010010" else
--"0000000010100000" when sig_inp <= "000000000000000000101010100011110101" else
--"0000000010011111" when sig_inp <= "000000000000000000101010100110000111" else
--"0000000010011110" when sig_inp <= "000000000000000000101010101000011001" else
--"0000000010011101" when sig_inp <= "000000000000000000101010101100111100" else
--"0000000010011100" when sig_inp <= "000000000000000000101010101111001101" else
--"0000000010011011" when sig_inp <= "000000000000000000101010110011110001" else
--"0000000010011010" when sig_inp <= "000000000000000000101010110110000010" else
--"0000000010011001" when sig_inp <= "000000000000000000101010111010100110" else
--"0000000010011000" when sig_inp <= "000000000000000000101010111100110111" else
--"0000000010010111" when sig_inp <= "000000000000000000101010111111001001" else
--"0000000010010110" when sig_inp <= "000000000000000000101011000011101100" else
--"0000000010010101" when sig_inp <= "000000000000000000101011000101111110" else
--"0000000010010100" when sig_inp <= "000000000000000000101011001010100001" else
--"0000000010010011" when sig_inp <= "000000000000000000101011001100110011" else
--"0000000010010010" when sig_inp <= "000000000000000000101011010001010110" else
--"0000000010010001" when sig_inp <= "000000000000000000101011010101111001" else
--"0000000010010000" when sig_inp <= "000000000000000000101011011000001011" else
--"0000000010001111" when sig_inp <= "000000000000000000101011011100101110" else
--"0000000010001110" when sig_inp <= "000000000000000000101011011111000000" else
--"0000000010001101" when sig_inp <= "000000000000000000101011100011100011" else
--"0000000010001100" when sig_inp <= "000000000000000000101011100101110101" else
--"0000000010001011" when sig_inp <= "000000000000000000101011101010011000" else
--"0000000010001010" when sig_inp <= "000000000000000000101011101110111011" else
--"0000000010001001" when sig_inp <= "000000000000000000101011110001001101" else
--"0000000010001000" when sig_inp <= "000000000000000000101011110101110000" else
--"0000000010000111" when sig_inp <= "000000000000000000101011111010010011" else
--"0000000010000110" when sig_inp <= "000000000000000000101011111100100101" else
--"0000000010000101" when sig_inp <= "000000000000000000101100000001001000" else
--"0000000010000100" when sig_inp <= "000000000000000000101100000101101100" else
--"0000000010000011" when sig_inp <= "000000000000000000101100000111111101" else
--"0000000010000010" when sig_inp <= "000000000000000000101100001100100000" else
--"0000000010000001" when sig_inp <= "000000000000000000101100010001000100" else
--"0000000010000000" when sig_inp <= "000000000000000000101100010011010101" else
--"0000000001111111" when sig_inp <= "000000000000000000101100010111111001" else
--"0000000001111110" when sig_inp <= "000000000000000000101100011100011100" else
--"0000000001111101" when sig_inp <= "000000000000000000101100100000111111" else
--"0000000001111100" when sig_inp <= "000000000000000000101100100101100010" else
--"0000000001111011" when sig_inp <= "000000000000000000101100100111110100" else
--"0000000001111010" when sig_inp <= "000000000000000000101100101100010111" else
--"0000000001111001" when sig_inp <= "000000000000000000101100110000111011" else
--"0000000001111000" when sig_inp <= "000000000000000000101100110101011110" else
--"0000000001110111" when sig_inp <= "000000000000000000101100111010000001" else
--"0000000001110110" when sig_inp <= "000000000000000000101100111110100100" else
--"0000000001110101" when sig_inp <= "000000000000000000101101000000110110" else
--"0000000001110100" when sig_inp <= "000000000000000000101101000101011001" else
--"0000000001110011" when sig_inp <= "000000000000000000101101001001111101" else
--"0000000001110010" when sig_inp <= "000000000000000000101101001110100000" else
--"0000000001110001" when sig_inp <= "000000000000000000101101010011000011" else
--"0000000001110000" when sig_inp <= "000000000000000000101101010111100110" else
--"0000000001101111" when sig_inp <= "000000000000000000101101011100001010" else
--"0000000001101110" when sig_inp <= "000000000000000000101101100000101101" else
--"0000000001101101" when sig_inp <= "000000000000000000101101100101010000" else
--"0000000001101100" when sig_inp <= "000000000000000000101101101001110100" else
--"0000000001101011" when sig_inp <= "000000000000000000101101101110010111" else
--"0000000001101010" when sig_inp <= "000000000000000000101101110010111010" else
--"0000000001101001" when sig_inp <= "000000000000000000101101111001101111" else
--"0000000001101000" when sig_inp <= "000000000000000000101101111110010010" else
--"0000000001100111" when sig_inp <= "000000000000000000101110000010110110" else
--"0000000001100110" when sig_inp <= "000000000000000000101110000111011001" else
--"0000000001100101" when sig_inp <= "000000000000000000101110001011111100" else
--"0000000001100100" when sig_inp <= "000000000000000000101110010000011111" else
--"0000000001100011" when sig_inp <= "000000000000000000101110010111010100" else
--"0000000001100010" when sig_inp <= "000000000000000000101110011011111000" else
--"0000000001100001" when sig_inp <= "000000000000000000101110100000011011" else
--"0000000001100000" when sig_inp <= "000000000000000000101110100111010000" else
--"0000000001011111" when sig_inp <= "000000000000000000101110101011110011" else
--"0000000001011110" when sig_inp <= "000000000000000000101110110000010110" else
--"0000000001011101" when sig_inp <= "000000000000000000101110110111001011" else
--"0000000001011100" when sig_inp <= "000000000000000000101110111011101110" else
--"0000000001011011" when sig_inp <= "000000000000000000101111000000010010" else
--"0000000001011010" when sig_inp <= "000000000000000000101111000111000111" else
--"0000000001011001" when sig_inp <= "000000000000000000101111001011101010" else
--"0000000001011000" when sig_inp <= "000000000000000000101111010010011111" else
--"0000000001010111" when sig_inp <= "000000000000000000101111010111000010" else
--"0000000001010110" when sig_inp <= "000000000000000000101111011101110111" else
--"0000000001010101" when sig_inp <= "000000000000000000101111100100101100" else
--"0000000001010100" when sig_inp <= "000000000000000000101111101001001111" else
--"0000000001010011" when sig_inp <= "000000000000000000101111110000000100" else
--"0000000001010010" when sig_inp <= "000000000000000000101111110110111001" else
--"0000000001010001" when sig_inp <= "000000000000000000101111111011011100" else
--"0000000001010000" when sig_inp <= "000000000000000000110000000010010001" else
--"0000000001001111" when sig_inp <= "000000000000000000110000001001000110" else
--"0000000001001110" when sig_inp <= "000000000000000000110000001111111011" else
--"0000000001001101" when sig_inp <= "000000000000000000110000010110110000" else
--"0000000001001100" when sig_inp <= "000000000000000000110000011101100101" else
--"0000000001001011" when sig_inp <= "000000000000000000110000100010001000" else
--"0000000001001010" when sig_inp <= "000000000000000000110000101000111101" else
--"0000000001001001" when sig_inp <= "000000000000000000110000101111110010" else
--"0000000001001000" when sig_inp <= "000000000000000000110000111000111000" else
--"0000000001000111" when sig_inp <= "000000000000000000110000111111101101" else
--"0000000001000110" when sig_inp <= "000000000000000000110001000110100010" else
--"0000000001000101" when sig_inp <= "000000000000000000110001001101010111" else
--"0000000001000100" when sig_inp <= "000000000000000000110001010100001100" else
--"0000000001000011" when sig_inp <= "000000000000000000110001011011000001" else
--"0000000001000010" when sig_inp <= "000000000000000000110001100100000111" else
--"0000000001000001" when sig_inp <= "000000000000000000110001101010111100" else
--"0000000001000000" when sig_inp <= "000000000000000000110001110100000011" else
--"0000000000111111" when sig_inp <= "000000000000000000110001111010111000" else
--"0000000000111110" when sig_inp <= "000000000000000000110010000011111110" else
--"0000000000111101" when sig_inp <= "000000000000000000110010001010110011" else
--"0000000000111100" when sig_inp <= "000000000000000000110010010011111010" else
--"0000000000111011" when sig_inp <= "000000000000000000110010011101000000" else
--"0000000000111010" when sig_inp <= "000000000000000000110010100011110101" else
--"0000000000111001" when sig_inp <= "000000000000000000110010101100111100" else
--"0000000000111000" when sig_inp <= "000000000000000000110010110110000010" else
--"0000000000110111" when sig_inp <= "000000000000000000110010111111001001" else
--"0000000000110110" when sig_inp <= "000000000000000000110011001000001111" else
--"0000000000110101" when sig_inp <= "000000000000000000110011010001010110" else
--"0000000000110100" when sig_inp <= "000000000000000000110011011100101110" else
--"0000000000110011" when sig_inp <= "000000000000000000110011100101110101" else
--"0000000000110010" when sig_inp <= "000000000000000000110011101110111011" else
--"0000000000110001" when sig_inp <= "000000000000000000110011111010010011" else
--"0000000000110000" when sig_inp <= "000000000000000000110100000011011010" else
--"0000000000101111" when sig_inp <= "000000000000000000110100001110110010" else
--"0000000000101110" when sig_inp <= "000000000000000000110100011010001010" else
--"0000000000101101" when sig_inp <= "000000000000000000110100100011010001" else
--"0000000000101100" when sig_inp <= "000000000000000000110100101110101001" else
--"0000000000101011" when sig_inp <= "000000000000000000110100111010000001" else
--"0000000000101010" when sig_inp <= "000000000000000000110101000111101011" else
--"0000000000101001" when sig_inp <= "000000000000000000110101010011000011" else
--"0000000000101000" when sig_inp <= "000000000000000000110101011110011011" else
--"0000000000100111" when sig_inp <= "000000000000000000110101101100000101" else
--"0000000000100110" when sig_inp <= "000000000000000000110101111001101111" else
--"0000000000100101" when sig_inp <= "000000000000000000110110000101000111" else
--"0000000000100100" when sig_inp <= "000000000000000000110110010010110001" else
--"0000000000100011" when sig_inp <= "000000000000000000110110100010101100" else
--"0000000000100010" when sig_inp <= "000000000000000000110110110000010110" else
--"0000000000100001" when sig_inp <= "000000000000000000110110111110000000" else
--"0000000000100000" when sig_inp <= "000000000000000000110111001101111100" else
--"0000000000011111" when sig_inp <= "000000000000000000110111011101110111" else
--"0000000000011110" when sig_inp <= "000000000000000000110111101101110010" else
--"0000000000011101" when sig_inp <= "000000000000000000111000000000000000" else
--"0000000000011100" when sig_inp <= "000000000000000000111000001111111011" else
--"0000000000011011" when sig_inp <= "000000000000000000111000100010001000" else
--"0000000000011010" when sig_inp <= "000000000000000000111000110100010101" else
--"0000000000011001" when sig_inp <= "000000000000000000111001001000110100" else
--"0000000000011000" when sig_inp <= "000000000000000000111001011101010011" else
--"0000000000010111" when sig_inp <= "000000000000000000111001110001110001" else
--"0000000000010110" when sig_inp <= "000000000000000000111010000110010000" else
--"0000000000010101" when sig_inp <= "000000000000000000111010011101000000" else
--"0000000000010100" when sig_inp <= "000000000000000000111010110110000010" else
--"0000000000010011" when sig_inp <= "000000000000000000111011001111000100" else
--"0000000000010010" when sig_inp <= "000000000000000000111011101000000110" else
--"0000000000010001" when sig_inp <= "000000000000000000111100000101101100" else
--"0000000000010000" when sig_inp <= "000000000000000000111100100000111111" else
--"0000000000001111" when sig_inp <= "000000000000000000111101000000110110" else
--"0000000000001110" when sig_inp <= "000000000000000000111101100010111111" else
--"0000000000001101" when sig_inp <= "000000000000000000111110000101000111" else
--"0000000000001100" when sig_inp <= "000000000000000000111110101011110011" else
--"0000000000001011" when sig_inp <= "000000000000000000111111010100110000" else
--"0000000000001010" when sig_inp <= "000000000000000001000000000000000000" else
--"0000000000001001" when sig_inp <= "000000000000000001000000110010000011" else
--"0000000000001000" when sig_inp <= "000000000000000001000001100110011001" else
--"0000000000000111" when sig_inp <= "000000000000000001000010100011110101" else
--"0000000000000110" when sig_inp <= "000000000000000001000011101000000110" else
--"0000000000000101" when sig_inp <= "000000000000000001000100110111110000" else
--"0000000000000100" when sig_inp <= "000000000000000001000110010101000011" else
--"0000000000000011" when sig_inp <= "000000000000000001001000000110110100" else
--"0000000000000010" when sig_inp <= "000000000000000001001010011010101111" else
--"0000000000000001" when sig_inp <= "000000000000000001001101101001110100" else
--"0000000000000000" when sig_inp <= "000000000000000001010011001100110011" else
--"0000000000000000";

--"1000000000000000" when sig_inp = "00000000000000000000" else
--"0111110101110111" when sig_inp <= "00000000001010001111" else
--"0111101011111011" when sig_inp <= "00000000010100011110" else
--"0111100010001011" when sig_inp <= "00000000011110101110" else
--"0111011000101000" when sig_inp <= "00000000101000111101" else
--"0111001111010001" when sig_inp <= "00000000110011001100" else
--"0111000110000110" when sig_inp <= "00000000111101011100" else
--"0110111101000111" when sig_inp <= "00000001000111101011" else
--"0110110100010011" when sig_inp <= "00000001010001111010" else
--"0110101011101010" when sig_inp <= "00000001011100001010" else
--"0110100011001100" when sig_inp <= "00000001100110011001" else
--"0110011010111000" when sig_inp <= "00000001110000101000" else
--"0110010010110000" when sig_inp <= "00000001111010111000" else
--"0110001010110001" when sig_inp <= "00000010000101000111" else
--"0110000010111101" when sig_inp <= "00000010001111010111" else
--"0101111011010011" when sig_inp <= "00000010011001100110" else
--"0101110011110010" when sig_inp <= "00000010100011110101" else
--"0101101100011011" when sig_inp <= "00000010101110000101" else
--"0101100101001101" when sig_inp <= "00000010111000010100" else
--"0101011110001000" when sig_inp <= "00000011000010100011" else
--"0101010111001101" when sig_inp <= "00000011001100110011" else
--"0101010000011010" when sig_inp <= "00000011010111000010" else
--"0101001001101111" when sig_inp <= "00000011100001010001" else
--"0101000011001101" when sig_inp <= "00000011101011100001" else
--"0100111100110100" when sig_inp <= "00000011110101110000" else
--"0100110110100010" when sig_inp <= "00000100000000000000" else
--"0100110000011001" when sig_inp <= "00000100001010001111" else
--"0100101010010111" when sig_inp <= "00000100010100011110" else
--"0100100100011101" when sig_inp <= "00000100011110101110" else
--"0100011110101010" when sig_inp <= "00000100101000111101" else
--"0100011000111111" when sig_inp <= "00000100110011001100" else
--"0100010011011011" when sig_inp <= "00000100111101011100" else
--"0100001101111110" when sig_inp <= "00000101000111101011" else
--"0100001000101000" when sig_inp <= "00000101010001111010" else
--"0100000011011000" when sig_inp <= "00000101011100001010" else
--"0011111110010000" when sig_inp <= "00000101100110011001" else
--"0011111001001101" when sig_inp <= "00000101110000101000" else
--"0011110100010010" when sig_inp <= "00000101111010111000" else
--"0011101111011100" when sig_inp <= "00000110000101000111" else
--"0011101010101101" when sig_inp <= "00000110001111010111" else
--"0011100110000011" when sig_inp <= "00000110011001100110" else
--"0011100001100000" when sig_inp <= "00000110100011110101" else
--"0011011101000010" when sig_inp <= "00000110101110000101" else
--"0011011000101010" when sig_inp <= "00000110111000010100" else
--"0011010100010111" when sig_inp <= "00000111000010100011" else
--"0011010000001010" when sig_inp <= "00000111001100110011" else
--"0011001100000010" when sig_inp <= "00000111010111000010" else
--"0011001000000000" when sig_inp <= "00000111100001010001" else
--"0011000100000010" when sig_inp <= "00000111101011100001" else
--"0011000000001010" when sig_inp <= "00000111110101110000" else
--"0010111100010110" when sig_inp <= "00001000000000000000" else
--"0010111000100111" when sig_inp <= "00001000001010001111" else
--"0010110100111110" when sig_inp <= "00001000010100011110" else
--"0010110001011000" when sig_inp <= "00001000011110101110" else
--"0010101101110111" when sig_inp <= "00001000101000111101" else
--"0010101010011011" when sig_inp <= "00001000110011001100" else
--"0010100111000011" when sig_inp <= "00001000111101011100" else
--"0010100011101111" when sig_inp <= "00001001000111101011" else
--"0010100000100000" when sig_inp <= "00001001010001111010" else
--"0010011101010100" when sig_inp <= "00001001011100001010" else
--"0010011010001101" when sig_inp <= "00001001100110011001" else
--"0010010111001010" when sig_inp <= "00001001110000101000" else
--"0010010100001010" when sig_inp <= "00001001111010111000" else
--"0010010001001110" when sig_inp <= "00001010000101000111" else
--"0010001110010110" when sig_inp <= "00001010001111010111" else
--"0010001011100010" when sig_inp <= "00001010011001100110" else
--"0010001000110001" when sig_inp <= "00001010100011110101" else
--"0010000110000100" when sig_inp <= "00001010101110000101" else
--"0010000011011010" when sig_inp <= "00001010111000010100" else
--"0010000000110011" when sig_inp <= "00001011000010100011" else
--"0001111110010000" when sig_inp <= "00001011001100110011" else
--"0001111011110000" when sig_inp <= "00001011010111000010" else
--"0001111001010011" when sig_inp <= "00001011100001010001" else
--"0001110110111001" when sig_inp <= "00001011101011100001" else
--"0001110100100011" when sig_inp <= "00001011110101110000" else
--"0001110010001111" when sig_inp <= "00001100000000000000" else
--"0001101111111110" when sig_inp <= "00001100001010001111" else
--"0001101101110000" when sig_inp <= "00001100010100011110" else
--"0001101011100101" when sig_inp <= "00001100011110101110" else
--"0001101001011101" when sig_inp <= "00001100101000111101" else
--"0001100111010111" when sig_inp <= "00001100110011001100" else
--"0001100101010100" when sig_inp <= "00001100111101011100" else
--"0001100011010100" when sig_inp <= "00001101000111101011" else
--"0001100001010110" when sig_inp <= "00001101010001111010" else
--"0001011111011011" when sig_inp <= "00001101011100001010" else
--"0001011101100010" when sig_inp <= "00001101100110011001" else
--"0001011011101011" when sig_inp <= "00001101110000101000" else
--"0001011001110111" when sig_inp <= "00001101111010111000" else
--"0001011000000101" when sig_inp <= "00001110000101000111" else
--"0001010110010101" when sig_inp <= "00001110001111010111" else
--"0001010100101000" when sig_inp <= "00001110011001100110" else
--"0001010010111101" when sig_inp <= "00001110100011110101" else
--"0001010001010100" when sig_inp <= "00001110101110000101" else
--"0001001111101101" when sig_inp <= "00001110111000010100" else
--"0001001110001000" when sig_inp <= "00001111000010100011" else
--"0001001100100101" when sig_inp <= "00001111001100110011" else
--"0001001011000100" when sig_inp <= "00001111010111000010" else
--"0001001001100100" when sig_inp <= "00001111100001010001" else
--"0001001000000111" when sig_inp <= "00001111101011100001" else
--"0001000110101100" when sig_inp <= "00001111110101110000" else
--"0001000101010010" when sig_inp <= "00010000000000000000" else
--"0001000011111010" when sig_inp <= "00010000001010001111" else
--"0001000010100100" when sig_inp <= "00010000010100011110" else
--"0001000001010000" when sig_inp <= "00010000011110101110" else
--"0000111111111101" when sig_inp <= "00010000101000111101" else
--"0000111110101100" when sig_inp <= "00010000110011001100" else
--"0000111101011101" when sig_inp <= "00010000111101011100" else
--"0000111100001111" when sig_inp <= "00010001000111101011" else
--"0000111011000010" when sig_inp <= "00010001010001111010" else
--"0000111001111000" when sig_inp <= "00010001011100001010" else
--"0000111000101110" when sig_inp <= "00010001100110011001" else
--"0000110111100110" when sig_inp <= "00010001110000101000" else
--"0000110110100000" when sig_inp <= "00010001111010111000" else
--"0000110101011011" when sig_inp <= "00010010000101000111" else
--"0000110100010111" when sig_inp <= "00010010001111010111" else
--"0000110011010101" when sig_inp <= "00010010011001100110" else
--"0000110010010100" when sig_inp <= "00010010100011110101" else
--"0000110001010100" when sig_inp <= "00010010101110000101" else
--"0000110000010101" when sig_inp <= "00010010111000010100" else
--"0000101111011000" when sig_inp <= "00010011000010100011" else
--"0000101110011100" when sig_inp <= "00010011001100110011" else
--"0000101101100001" when sig_inp <= "00010011010111000010" else
--"0000101100101000" when sig_inp <= "00010011100001010001" else
--"0000101011101111" when sig_inp <= "00010011101011100001" else
--"0000101010111000" when sig_inp <= "00010011110101110000" else
--"0000101010000001" when sig_inp <= "00010100000000000000" else
--"0000101001001100" when sig_inp <= "00010100001010001111" else
--"0000101000011000" when sig_inp <= "00010100010100011110" else
--"0000100111100101" when sig_inp <= "00010100011110101110" else
--"0000100110110010" when sig_inp <= "00010100101000111101" else
--"0000100110000001" when sig_inp <= "00010100110011001100" else
--"0000100101010001" when sig_inp <= "00010100111101011100" else
--"0000100100100010" when sig_inp <= "00010101000111101011" else
--"0000100011110100" when sig_inp <= "00010101010001111010" else
--"0000100011000110" when sig_inp <= "00010101011100001010" else
--"0000100010011010" when sig_inp <= "00010101100110011001" else
--"0000100001101110" when sig_inp <= "00010101110000101000" else
--"0000100001000011" when sig_inp <= "00010101111010111000" else
--"0000100000011001" when sig_inp <= "00010110000101000111" else
--"0000011111110000" when sig_inp <= "00010110001111010111" else
--"0000011111001000" when sig_inp <= "00010110011001100110" else
--"0000011110100001" when sig_inp <= "00010110100011110101" else
--"0000011101111010" when sig_inp <= "00010110101110000101" else
--"0000011101010100" when sig_inp <= "00010110111000010100" else
--"0000011100101111" when sig_inp <= "00010111000010100011" else
--"0000011100001011" when sig_inp <= "00010111001100110011" else
--"0000011011100111" when sig_inp <= "00010111010111000010" else
--"0000011011000100" when sig_inp <= "00010111100001010001" else
--"0000011010100010" when sig_inp <= "00010111101011100001" else
--"0000011010000000" when sig_inp <= "00010111110101110000" else
--"0000011001011111" when sig_inp <= "00011000000000000000" else
--"0000011000111111" when sig_inp <= "00011000001010001111" else
--"0000011000011111" when sig_inp <= "00011000010100011110" else
--"0000011000000000" when sig_inp <= "00011000011110101110" else
--"0000010111100001" when sig_inp <= "00011000101000111101" else
--"0000010111000100" when sig_inp <= "00011000110011001100" else
--"0000010110100110" when sig_inp <= "00011000111101011100" else
--"0000010110001010" when sig_inp <= "00011001000111101011" else
--"0000010101101110" when sig_inp <= "00011001010001111010" else
--"0000010101010010" when sig_inp <= "00011001011100001010" else
--"0000010100110111" when sig_inp <= "00011001100110011001" else
--"0000010100011101" when sig_inp <= "00011001110000101000" else
--"0000010100000011" when sig_inp <= "00011001111010111000" else
--"0000010011101001" when sig_inp <= "00011010000101000111" else
--"0000010011010001" when sig_inp <= "00011010001111010111" else
--"0000010010111000" when sig_inp <= "00011010011001100110" else
--"0000010010100000" when sig_inp <= "00011010100011110101" else
--"0000010010001001" when sig_inp <= "00011010101110000101" else
--"0000010001110010" when sig_inp <= "00011010111000010100" else
--"0000010001011011" when sig_inp <= "00011011000010100011" else
--"0000010001000101" when sig_inp <= "00011011001100110011" else
--"0000010000101111" when sig_inp <= "00011011010111000010" else
--"0000010000011010" when sig_inp <= "00011011100001010001" else
--"0000010000000101" when sig_inp <= "00011011101011100001" else
--"0000001111110001" when sig_inp <= "00011011110101110000" else
--"0000001111011101" when sig_inp <= "00011100000000000000" else
--"0000001111001001" when sig_inp <= "00011100001010001111" else
--"0000001110110110" when sig_inp <= "00011100010100011110" else
--"0000001110100011" when sig_inp <= "00011100011110101110" else
--"0000001110010001" when sig_inp <= "00011100101000111101" else
--"0000001101111111" when sig_inp <= "00011100110011001100" else
--"0000001101101101" when sig_inp <= "00011100111101011100" else
--"0000001101011100" when sig_inp <= "00011101000111101011" else
--"0000001101001011" when sig_inp <= "00011101010001111010" else
--"0000001100111010" when sig_inp <= "00011101011100001010" else
--"0000001100101010" when sig_inp <= "00011101100110011001" else
--"0000001100011010" when sig_inp <= "00011101110000101000" else
--"0000001100001010" when sig_inp <= "00011101111010111000" else
--"0000001011111010" when sig_inp <= "00011110000101000111" else
--"0000001011101011" when sig_inp <= "00011110001111010111" else
--"0000001011011101" when sig_inp <= "00011110011001100110" else
--"0000001011001110" when sig_inp <= "00011110100011110101" else
--"0000001011000000" when sig_inp <= "00011110101110000101" else
--"0000001010110010" when sig_inp <= "00011110111000010100" else
--"0000001010100100" when sig_inp <= "00011111000010100011" else
--"0000001010010111" when sig_inp <= "00011111001100110011" else
--"0000001010001010" when sig_inp <= "00011111010111000010" else
--"0000001001111101" when sig_inp <= "00011111100001010001" else
--"0000001001110000" when sig_inp <= "00011111101011100001" else
--"0000001001100100" when sig_inp <= "00011111110101110000" else
--"0000001001011000" when sig_inp <= "00100000000000000000" else
--"0000001001001100" when sig_inp <= "00100000001010001111" else
--"0000001001000000" when sig_inp <= "00100000010100011110" else
--"0000001000110101" when sig_inp <= "00100000011110101110" else
--"0000001000101010" when sig_inp <= "00100000101000111101" else
--"0000001000011111" when sig_inp <= "00100000110011001100" else
--"0000001000010100" when sig_inp <= "00100000111101011100" else
--"0000001000001001" when sig_inp <= "00100001000111101011" else
--"0000000111111111" when sig_inp <= "00100001010001111010" else
--"0000000111110101" when sig_inp <= "00100001011100001010" else
--"0000000111101011" when sig_inp <= "00100001100110011001" else
--"0000000111100001" when sig_inp <= "00100001110000101000" else
--"0000000111011000" when sig_inp <= "00100001111010111000" else
--"0000000111001110" when sig_inp <= "00100010000101000111" else
--"0000000111000101" when sig_inp <= "00100010001111010111" else
--"0000000110111100" when sig_inp <= "00100010011001100110" else
--"0000000110110011" when sig_inp <= "00100010100011110101" else
--"0000000110101011" when sig_inp <= "00100010101110000101" else
--"0000000110100010" when sig_inp <= "00100010111000010100" else
--"0000000110011010" when sig_inp <= "00100011000010100011" else
--"0000000110010010" when sig_inp <= "00100011001100110011" else
--"0000000110001010" when sig_inp <= "00100011010111000010" else
--"0000000110000010" when sig_inp <= "00100011100001010001" else
--"0000000101111010" when sig_inp <= "00100011101011100001" else
--"0000000101110011" when sig_inp <= "00100011110101110000" else
--"0000000101101100" when sig_inp <= "00100100000000000000" else
--"0000000101100100" when sig_inp <= "00100100001010001111" else
--"0000000101011101" when sig_inp <= "00100100010100011110" else
--"0000000101010110" when sig_inp <= "00100100011110101110" else
--"0000000101010000" when sig_inp <= "00100100101000111101" else
--"0000000101001001" when sig_inp <= "00100100110011001100" else
--"0000000101000010" when sig_inp <= "00100100111101011100" else
--"0000000100111100" when sig_inp <= "00100101000111101011" else
--"0000000100110110" when sig_inp <= "00100101010001111010" else
--"0000000100110000" when sig_inp <= "00100101011100001010" else
--"0000000100101010" when sig_inp <= "00100101100110011001" else
--"0000000100100100" when sig_inp <= "00100101110000101000" else
--"0000000100011110" when sig_inp <= "00100101111010111000" else
--"0000000100011000" when sig_inp <= "00100110000101000111" else
--"0000000100010011" when sig_inp <= "00100110001111010111" else
--"0000000100001101" when sig_inp <= "00100110011001100110" else
--"0000000100001000" when sig_inp <= "00100110100011110101" else
--"0000000100000011" when sig_inp <= "00100110101110000101" else
--"0000000011111101" when sig_inp <= "00100110111000010100" else
--"0000000011111000" when sig_inp <= "00100111000010100011" else
--"0000000011110100" when sig_inp <= "00100111001100110011" else
--"0000000011101111" when sig_inp <= "00100111010111000010" else
--"0000000011101010" when sig_inp <= "00100111100001010001" else
--"0000000011100101" when sig_inp <= "00100111101011100001" else
--"0000000011100001" when sig_inp <= "00100111110101110000" else
--"0000000011011100" when sig_inp <= "00101000000000000000" else
--"0000000011011000" when sig_inp <= "00101000001010001111" else
--"0000000011010100" when sig_inp <= "00101000010100011110" else
--"0000000011001111" when sig_inp <= "00101000011110101110" else
--"0000000011001011" when sig_inp <= "00101000101000111101" else
--"0000000011000111" when sig_inp <= "00101000110011001100" else
--"0000000011000011" when sig_inp <= "00101000111101011100" else
--"0000000010111111" when sig_inp <= "00101001000111101011" else
--"0000000010111100" when sig_inp <= "00101001010001111010" else
--"0000000010111000" when sig_inp <= "00101001011100001010" else
--"0000000010110100" when sig_inp <= "00101001100110011001" else
--"0000000010110001" when sig_inp <= "00101001110000101000" else
--"0000000010101101" when sig_inp <= "00101001111010111000" else
--"0000000010101010" when sig_inp <= "00101010000101000111" else
--"0000000010100110" when sig_inp <= "00101010001111010111" else
--"0000000010100011" when sig_inp <= "00101010011001100110" else
--"0000000010100000" when sig_inp <= "00101010100011110101" else
--"0000000010011101" when sig_inp <= "00101010101110000101" else
--"0000000010011010" when sig_inp <= "00101010111000010100" else
--"0000000010010110" when sig_inp <= "00101011000010100011" else
--"0000000010010011" when sig_inp <= "00101011001100110011" else
--"0000000010010001" when sig_inp <= "00101011010111000010" else
--"0000000010001110" when sig_inp <= "00101011100001010001" else
--"0000000010001011" when sig_inp <= "00101011101011100001" else
--"0000000010001000" when sig_inp <= "00101011110101110000" else
--"0000000010000101" when sig_inp <= "00101100000000000000" else
--"0000000010000011" when sig_inp <= "00101100001010001111" else
--"0000000010000000" when sig_inp <= "00101100010100011110" else
--"0000000001111110" when sig_inp <= "00101100011110101110" else
--"0000000001111011" when sig_inp <= "00101100101000111101" else
--"0000000001111001" when sig_inp <= "00101100110011001100" else
--"0000000001110110" when sig_inp <= "00101100111101011100" else
--"0000000001110100" when sig_inp <= "00101101000111101011" else
--"0000000001110010" when sig_inp <= "00101101010001111010" else
--"0000000001101111" when sig_inp <= "00101101011100001010" else
--"0000000001101101" when sig_inp <= "00101101100110011001" else
--"0000000001101011" when sig_inp <= "00101101110000101000" else
--"0000000001101001" when sig_inp <= "00101101111010111000" else
--"0000000001100111" when sig_inp <= "00101110000101000111" else
--"0000000001100101" when sig_inp <= "00101110001111010111" else
--"0000000001100011" when sig_inp <= "00101110011001100110" else
--"0000000001100001" when sig_inp <= "00101110100011110101" else
--"0000000001011111" when sig_inp <= "00101110101110000101" else
--"0000000001011101" when sig_inp <= "00101110111000010100" else
--"0000000001011011" when sig_inp <= "00101111000010100011" else
--"0000000001011001" when sig_inp <= "00101111001100110011" else
--"0000000001010111" when sig_inp <= "00101111010111000010" else
--"0000000001010110" when sig_inp <= "00101111100001010001" else
--"0000000001010100" when sig_inp <= "00101111101011100001" else
--"0000000001010010" when sig_inp <= "00101111110101110000" else
--"0000000001010001" when sig_inp <= "00110000000000000000" else
--"0000000001001111" when sig_inp <= "00110000001010001111" else
--"0000000001001110" when sig_inp <= "00110000010100011110" else
--"0000000001001100" when sig_inp <= "00110000011110101110" else
--"0000000001001010" when sig_inp <= "00110000101000111101" else
--"0000000001001001" when sig_inp <= "00110000110011001100" else
--"0000000001001000" when sig_inp <= "00110000111101011100" else
--"0000000001000110" when sig_inp <= "00110001000111101011" else
--"0000000001000101" when sig_inp <= "00110001010001111010" else
--"0000000001000011" when sig_inp <= "00110001011100001010" else
--"0000000001000010" when sig_inp <= "00110001100110011001" else
--"0000000001000001" when sig_inp <= "00110001110000101000" else
--"0000000000111111" when sig_inp <= "00110001111010111000" else
--"0000000000111110" when sig_inp <= "00110010000101000111" else
--"0000000000111101" when sig_inp <= "00110010001111010111" else
--"0000000000111100" when sig_inp <= "00110010011001100110" else
--"0000000000111010" when sig_inp <= "00110010100011110101" else
--"0000000000111001" when sig_inp <= "00110010101110000101" else
--"0000000000111000" when sig_inp <= "00110010111000010100" else
--"0000000000110111" when sig_inp <= "00110011000010100011" else
--"0000000000110110" when sig_inp <= "00110011001100110011" else
--"0000000000110101" when sig_inp <= "00110011010111000010" else
--"0000000000110100" when sig_inp <= "00110011100001010001" else
--"0000000000110011" when sig_inp <= "00110011101011100001" else
--"0000000000110010" when sig_inp <= "00110011110101110000" else
--"0000000000110001" when sig_inp <= "00110100000000000000" else
--"0000000000110000" when sig_inp <= "00110100001010001111" else
--"0000000000101111" when sig_inp <= "00110100010100011110" else
--"0000000000101110" when sig_inp <= "00110100011110101110" else
--"0000000000101101" when sig_inp <= "00110100101000111101" else
--"0000000000101100" when sig_inp <= "00110100110011001100" else
--"0000000000101011" when sig_inp <= "00110100111101011100" else
--"0000000000101010" when sig_inp <= "00110101000111101011" else
--"0000000000101001" when sig_inp <= "00110101010001111010" else
--"0000000000101000" when sig_inp <= "00110101100110011001" else
--"0000000000100111" when sig_inp <= "00110101110000101000" else
--"0000000000100110" when sig_inp <= "00110101111010111000" else
--"0000000000100101" when sig_inp <= "00110110000101000111" else
--"0000000000100100" when sig_inp <= "00110110011001100110" else
--"0000000000100011" when sig_inp <= "00110110100011110101" else
--"0000000000100010" when sig_inp <= "00110110111000010100" else
--"0000000000100001" when sig_inp <= "00110111000010100011" else
--"0000000000100000" when sig_inp <= "00110111010111000010" else
--"0000000000011111" when sig_inp <= "00110111100001010001" else
--"0000000000011110" when sig_inp <= "00110111110101110000" else
--"0000000000011101" when sig_inp <= "00111000000000000000" else
--"0000000000011100" when sig_inp <= "00111000010100011110" else
--"0000000000011011" when sig_inp <= "00111000101000111101" else
--"0000000000011010" when sig_inp <= "00111000111101011100" else
--"0000000000011001" when sig_inp <= "00111001000111101011" else
--"0000000000011000" when sig_inp <= "00111001011100001010" else
--"0000000000010111" when sig_inp <= "00111001110000101000" else
--"0000000000010110" when sig_inp <= "00111010001111010111" else
--"0000000000010101" when sig_inp <= "00111010100011110101" else
--"0000000000010100" when sig_inp <= "00111010111000010100" else
--"0000000000010011" when sig_inp <= "00111011010111000010" else
--"0000000000010010" when sig_inp <= "00111011101011100001" else
--"0000000000010001" when sig_inp <= "00111100001010001111" else
--"0000000000010000" when sig_inp <= "00111100101000111101" else
--"0000000000001111" when sig_inp <= "00111101000111101011" else
--"0000000000001110" when sig_inp <= "00111101100110011001" else
--"0000000000001101" when sig_inp <= "00111110000101000111" else
--"0000000000001100" when sig_inp <= "00111110101110000101" else
--"0000000000001011" when sig_inp <= "00111111010111000010" else
--"0000000000001010" when sig_inp <= "01000000000000000000" else
--"0000000000001001" when sig_inp <= "01000000110011001100" else
--"0000000000001000" when sig_inp <= "01000001100110011001" else
--"0000000000000111" when sig_inp <= "01000010100011110101" else
--"0000000000000110" when sig_inp <= "01000011101011100001" else
--"0000000000000101" when sig_inp <= "01000100111101011100" else
--"0000000000000100" when sig_inp <= "01000110011001100110" else
--"0000000000000011" when sig_inp <= "01001000001010001111" else
--"0000000000000010" when sig_inp <= "01001010011001100110" else
--"0000000000000001" when sig_inp <= "01001101110000101000" else
--"0000000000000000";
----------------------------------------------------------------------------------------------------------------------------------------------------------------

--sig_out <= "1000000000000000" when sig_inp = "00000000000000000000" else
--"0111110101110111" when sig_inp <= "00000000001010001111" else
--"0111101011111011" when sig_inp <= "00000000010100011110" else
--"0111100010001011" when sig_inp <= "00000000011110101110" else
--"0111011000101000" when sig_inp <= "00000000101000111101" else
--"0111001111010001" when sig_inp <= "00000000110011001100" else
--"0111000110000110" when sig_inp <= "00000000111101011100" else
--"0110111101000111" when sig_inp <= "00000001000111101011" else
--"0110110100010011" when sig_inp <= "00000001010001111010" else
--"0110101011101010" when sig_inp <= "00000001011100001010" else
--"0110100011001100" when sig_inp <= "00000001100110011001" else
--"0110011010111000" when sig_inp <= "00000001110000101000" else
--"0110010010110000" when sig_inp <= "00000001111010111000" else
--"0110001010110001" when sig_inp <= "00000010000101000111" else
--"0110000010111101" when sig_inp <= "00000010001111010111" else
--"0101111011010011" when sig_inp <= "00000010011001100110" else
--"0101110011110010" when sig_inp <= "00000010100011110101" else
--"0101101100011011" when sig_inp <= "00000010101110000101" else
--"0101100101001101" when sig_inp <= "00000010111000010100" else
--"0101011110001000" when sig_inp <= "00000011000010100011" else
--"0101010111001101" when sig_inp <= "00000011001100110011" else
--"0101010000011010" when sig_inp <= "00000011010111000010" else
--"0101001001101111" when sig_inp <= "00000011100001010001" else
--"0101000011001101" when sig_inp <= "00000011101011100001" else
--"0100111100110100" when sig_inp <= "00000011110101110000" else
--"0100110110100010" when sig_inp <= "00000100000000000000" else
--"0100110000011001" when sig_inp <= "00000100001010001111" else
--"0100101010010111" when sig_inp <= "00000100010100011110" else
--"0100100100011101" when sig_inp <= "00000100011110101110" else
--"0100011110101010" when sig_inp <= "00000100101000111101" else
--"0100011000111111" when sig_inp <= "00000100110011001100" else
--"0100010011011011" when sig_inp <= "00000100111101011100" else
--"0100001101111110" when sig_inp <= "00000101000111101011" else
--"0100001000101000" when sig_inp <= "00000101010001111010" else
--"0100000011011000" when sig_inp <= "00000101011100001010" else
--"0011111110010000" when sig_inp <= "00000101100110011001" else
--"0011111001001101" when sig_inp <= "00000101110000101000" else
--"0011110100010010" when sig_inp <= "00000101111010111000" else
--"0011101111011100" when sig_inp <= "00000110000101000111" else
--"0011101010101101" when sig_inp <= "00000110001111010111" else
--"0011100110000011" when sig_inp <= "00000110011001100110" else
--"0011100001100000" when sig_inp <= "00000110100011110101" else
--"0011011101000010" when sig_inp <= "00000110101110000101" else
--"0011011000101010" when sig_inp <= "00000110111000010100" else
--"0011010100010111" when sig_inp <= "00000111000010100011" else
--"0011010000001010" when sig_inp <= "00000111001100110011" else
--"0011001100000010" when sig_inp <= "00000111010111000010" else
--"0011001000000000" when sig_inp <= "00000111100001010001" else
--"0011000100000010" when sig_inp <= "00000111101011100001" else
--"0011000000001010" when sig_inp <= "00000111110101110000" else
--"0010111100010110" when sig_inp <= "00001000000000000000" else
--"0010111000100111" when sig_inp <= "00001000001010001111" else
--"0010110100111110" when sig_inp <= "00001000010100011110" else
--"0010110001011000" when sig_inp <= "00001000011110101110" else
--"0010101101110111" when sig_inp <= "00001000101000111101" else
--"0010101010011011" when sig_inp <= "00001000110011001100" else
--"0010100111000011" when sig_inp <= "00001000111101011100" else
--"0010100011101111" when sig_inp <= "00001001000111101011" else
--"0010100000100000" when sig_inp <= "00001001010001111010" else
--"0010011101010100" when sig_inp <= "00001001011100001010" else
--"0010011010001101" when sig_inp <= "00001001100110011001" else
--"0010010111001010" when sig_inp <= "00001001110000101000" else
--"0010010100001010" when sig_inp <= "00001001111010111000" else
--"0010010001001110" when sig_inp <= "00001010000101000111" else
--"0010001110010110" when sig_inp <= "00001010001111010111" else
--"0010001011100010" when sig_inp <= "00001010011001100110" else
--"0010001000110001" when sig_inp <= "00001010100011110101" else
--"0010000110000100" when sig_inp <= "00001010101110000101" else
--"0010000011011010" when sig_inp <= "00001010111000010100" else
--"0010000000110011" when sig_inp <= "00001011000010100011" else
--"0001111110010000" when sig_inp <= "00001011001100110011" else
--"0001111011110000" when sig_inp <= "00001011010111000010" else
--"0001111001010011" when sig_inp <= "00001011100001010001" else
--"0001110110111001" when sig_inp <= "00001011101011100001" else
--"0001110100100011" when sig_inp <= "00001011110101110000" else
--"0001110010001111" when sig_inp <= "00001100000000000000" else
--"0001101111111110" when sig_inp <= "00001100001010001111" else
--"0001101101110000" when sig_inp <= "00001100010100011110" else
--"0001101011100101" when sig_inp <= "00001100011110101110" else
--"0001101001011101" when sig_inp <= "00001100101000111101" else
--"0001100111010111" when sig_inp <= "00001100110011001100" else
--"0001100101010100" when sig_inp <= "00001100111101011100" else
--"0001100011010100" when sig_inp <= "00001101000111101011" else
--"0001100001010110" when sig_inp <= "00001101010001111010" else
--"0001011111011011" when sig_inp <= "00001101011100001010" else
--"0001011101100010" when sig_inp <= "00001101100110011001" else
--"0001011011101011" when sig_inp <= "00001101110000101000" else
--"0001011001110111" when sig_inp <= "00001101111010111000" else
--"0001011000000101" when sig_inp <= "00001110000101000111" else
--"0001010110010101" when sig_inp <= "00001110001111010111" else
--"0001010100101000" when sig_inp <= "00001110011001100110" else
--"0001010010111101" when sig_inp <= "00001110100011110101" else
--"0001010001010100" when sig_inp <= "00001110101110000101" else
--"0001001111101101" when sig_inp <= "00001110111000010100" else
--"0001001110001000" when sig_inp <= "00001111000010100011" else
--"0001001100100101" when sig_inp <= "00001111001100110011" else
--"0001001011000100" when sig_inp <= "00001111010111000010" else
--"0001001001100100" when sig_inp <= "00001111100001010001" else
--"0001001000000111" when sig_inp <= "00001111101011100001" else
--"0001000110101100" when sig_inp <= "00001111110101110000" else
--"0001000101010010" when sig_inp <= "00010000000000000000" else
--"0001000011111010" when sig_inp <= "00010000001010001111" else
--"0001000010100100" when sig_inp <= "00010000010100011110" else
--"0001000001010000" when sig_inp <= "00010000011110101110" else
--"0000111111111101" when sig_inp <= "00010000101000111101" else
--"0000111110101100" when sig_inp <= "00010000110011001100" else
--"0000111101011101" when sig_inp <= "00010000111101011100" else
--"0000111100001111" when sig_inp <= "00010001000111101011" else
--"0000111011000010" when sig_inp <= "00010001010001111010" else
--"0000111001111000" when sig_inp <= "00010001011100001010" else
--"0000111000101110" when sig_inp <= "00010001100110011001" else
--"0000110111100110" when sig_inp <= "00010001110000101000" else
--"0000110110100000" when sig_inp <= "00010001111010111000" else
--"0000110101011011" when sig_inp <= "00010010000101000111" else
--"0000110100010111" when sig_inp <= "00010010001111010111" else
--"0000110011010101" when sig_inp <= "00010010011001100110" else
--"0000110010010100" when sig_inp <= "00010010100011110101" else
--"0000110001010100" when sig_inp <= "00010010101110000101" else
--"0000110000010101" when sig_inp <= "00010010111000010100" else
--"0000101111011000" when sig_inp <= "00010011000010100011" else
--"0000101110011100" when sig_inp <= "00010011001100110011" else
--"0000101101100001" when sig_inp <= "00010011010111000010" else
--"0000101100101000" when sig_inp <= "00010011100001010001" else
--"0000101011101111" when sig_inp <= "00010011101011100001" else
--"0000101010111000" when sig_inp <= "00010011110101110000" else
--"0000101010000001" when sig_inp <= "00010100000000000000" else
--"0000101001001100" when sig_inp <= "00010100001010001111" else
--"0000101000011000" when sig_inp <= "00010100010100011110" else
--"0000100111100101" when sig_inp <= "00010100011110101110" else
--"0000100110110010" when sig_inp <= "00010100101000111101" else
--"0000100110000001" when sig_inp <= "00010100110011001100" else
--"0000100101010001" when sig_inp <= "00010100111101011100" else
--"0000100100100010" when sig_inp <= "00010101000111101011" else
--"0000100011110100" when sig_inp <= "00010101010001111010" else
--"0000100011000110" when sig_inp <= "00010101011100001010" else
--"0000100010011010" when sig_inp <= "00010101100110011001" else
--"0000100001101110" when sig_inp <= "00010101110000101000" else
--"0000100001000011" when sig_inp <= "00010101111010111000" else
--"0000100000011001" when sig_inp <= "00010110000101000111" else
--"0000011111110000" when sig_inp <= "00010110001111010111" else
--"0000011111001000" when sig_inp <= "00010110011001100110" else
--"0000011110100001" when sig_inp <= "00010110100011110101" else
--"0000011101111010" when sig_inp <= "00010110101110000101" else
--"0000011101010100" when sig_inp <= "00010110111000010100" else
--"0000011100101111" when sig_inp <= "00010111000010100011" else
--"0000011100001011" when sig_inp <= "00010111001100110011" else
--"0000011011100111" when sig_inp <= "00010111010111000010" else
--"0000011011000100" when sig_inp <= "00010111100001010001" else
--"0000011010100010" when sig_inp <= "00010111101011100001" else
--"0000011010000000" when sig_inp <= "00010111110101110000" else
--"0000011001011111" when sig_inp <= "00011000000000000000" else
--"0000011000111111" when sig_inp <= "00011000001010001111" else
--"0000011000011111" when sig_inp <= "00011000010100011110" else
--"0000011000000000" when sig_inp <= "00011000011110101110" else
--"0000010111100001" when sig_inp <= "00011000101000111101" else
--"0000010111000100" when sig_inp <= "00011000110011001100" else
--"0000010110100110" when sig_inp <= "00011000111101011100" else
--"0000010110001010" when sig_inp <= "00011001000111101011" else
--"0000010101101110" when sig_inp <= "00011001010001111010" else
--"0000010101010010" when sig_inp <= "00011001011100001010" else
--"0000010100110111" when sig_inp <= "00011001100110011001" else
--"0000010100011101" when sig_inp <= "00011001110000101000" else
--"0000010100000011" when sig_inp <= "00011001111010111000" else
--"0000010011101001" when sig_inp <= "00011010000101000111" else
--"0000010011010001" when sig_inp <= "00011010001111010111" else
--"0000010010111000" when sig_inp <= "00011010011001100110" else
--"0000010010100000" when sig_inp <= "00011010100011110101" else
--"0000010010001001" when sig_inp <= "00011010101110000101" else
--"0000010001110010" when sig_inp <= "00011010111000010100" else
--"0000010001011011" when sig_inp <= "00011011000010100011" else
--"0000010001000101" when sig_inp <= "00011011001100110011" else
--"0000010000101111" when sig_inp <= "00011011010111000010" else
--"0000010000011010" when sig_inp <= "00011011100001010001" else
--"0000010000000101" when sig_inp <= "00011011101011100001" else
--"0000001111110001" when sig_inp <= "00011011110101110000" else
--"0000001111011101" when sig_inp <= "00011100000000000000" else
--"0000001111001001" when sig_inp <= "00011100001010001111" else
--"0000001110110110" when sig_inp <= "00011100010100011110" else
--"0000001110100011" when sig_inp <= "00011100011110101110" else
--"0000001110010001" when sig_inp <= "00011100101000111101" else
--"0000001101111111" when sig_inp <= "00011100110011001100" else
--"0000001101101101" when sig_inp <= "00011100111101011100" else
--"0000001101011100" when sig_inp <= "00011101000111101011" else
--"0000001101001011" when sig_inp <= "00011101010001111010" else
--"0000001100111010" when sig_inp <= "00011101011100001010" else
--"0000001100101010" when sig_inp <= "00011101100110011001" else
--"0000001100011010" when sig_inp <= "00011101110000101000" else
--"0000001100001010" when sig_inp <= "00011101111010111000" else
--"0000001011111010" when sig_inp <= "00011110000101000111" else
--"0000001011101011" when sig_inp <= "00011110001111010111" else
--"0000001011011101" when sig_inp <= "00011110011001100110" else
--"0000001011001110" when sig_inp <= "00011110100011110101" else
--"0000001011000000" when sig_inp <= "00011110101110000101" else
--"0000001010110010" when sig_inp <= "00011110111000010100" else
--"0000001010100100" when sig_inp <= "00011111000010100011" else
--"0000001010010111" when sig_inp <= "00011111001100110011" else
--"0000001010001010" when sig_inp <= "00011111010111000010" else
--"0000001001111101" when sig_inp <= "00011111100001010001" else
--"0000001001110000" when sig_inp <= "00011111101011100001" else
--"0000001001100100" when sig_inp <= "00011111110101110000" else
--"0000001001011000" when sig_inp <= "00100000000000000000" else
--"0000001001001100" when sig_inp <= "00100000001010001111" else
--"0000001001000000" when sig_inp <= "00100000010100011110" else
--"0000001000110101" when sig_inp <= "00100000011110101110" else
--"0000001000101010" when sig_inp <= "00100000101000111101" else
--"0000001000011111" when sig_inp <= "00100000110011001100" else
--"0000001000010100" when sig_inp <= "00100000111101011100" else
--"0000001000001001" when sig_inp <= "00100001000111101011" else
--"0000000111111111" when sig_inp <= "00100001010001111010" else
--"0000000111110101" when sig_inp <= "00100001011100001010" else
--"0000000111101011" when sig_inp <= "00100001100110011001" else
--"0000000111100001" when sig_inp <= "00100001110000101000" else
--"0000000111011000" when sig_inp <= "00100001111010111000" else
--"0000000111001110" when sig_inp <= "00100010000101000111" else
--"0000000111000101" when sig_inp <= "00100010001111010111" else
--"0000000110111100" when sig_inp <= "00100010011001100110" else
--"0000000110110011" when sig_inp <= "00100010100011110101" else
--"0000000110101011" when sig_inp <= "00100010101110000101" else
--"0000000110100010" when sig_inp <= "00100010111000010100" else
--"0000000110011010" when sig_inp <= "00100011000010100011" else
--"0000000110010010" when sig_inp <= "00100011001100110011" else
--"0000000110001010" when sig_inp <= "00100011010111000010" else
--"0000000110000010" when sig_inp <= "00100011100001010001" else
--"0000000101111010" when sig_inp <= "00100011101011100001" else
--"0000000101110011" when sig_inp <= "00100011110101110000" else
--"0000000101101100" when sig_inp <= "00100100000000000000" else
--"0000000101100100" when sig_inp <= "00100100001010001111" else
--"0000000101011101" when sig_inp <= "00100100010100011110" else
--"0000000101010110" when sig_inp <= "00100100011110101110" else
--"0000000101010000" when sig_inp <= "00100100101000111101" else
--"0000000101001001" when sig_inp <= "00100100110011001100" else
--"0000000101000010" when sig_inp <= "00100100111101011100" else
--"0000000100111100" when sig_inp <= "00100101000111101011" else
--"0000000100110110" when sig_inp <= "00100101010001111010" else
--"0000000100110000" when sig_inp <= "00100101011100001010" else
--"0000000100101010" when sig_inp <= "00100101100110011001" else
--"0000000100100100" when sig_inp <= "00100101110000101000" else
--"0000000100011110" when sig_inp <= "00100101111010111000" else
--"0000000100011000" when sig_inp <= "00100110000101000111" else
--"0000000100010011" when sig_inp <= "00100110001111010111" else
--"0000000100001101" when sig_inp <= "00100110011001100110" else
--"0000000100001000" when sig_inp <= "00100110100011110101" else
--"0000000100000011" when sig_inp <= "00100110101110000101" else
--"0000000011111101" when sig_inp <= "00100110111000010100" else
--"0000000011111000" when sig_inp <= "00100111000010100011" else
--"0000000011110100" when sig_inp <= "00100111001100110011" else
--"0000000011101111" when sig_inp <= "00100111010111000010" else
--"0000000011101010" when sig_inp <= "00100111100001010001" else
--"0000000011100101" when sig_inp <= "00100111101011100001" else
--"0000000011100001" when sig_inp <= "00100111110101110000" else
--"0000000011011100" when sig_inp <= "00101000000000000000" else
--"0000000011011000" when sig_inp <= "00101000001010001111" else
--"0000000011010100" when sig_inp <= "00101000010100011110" else
--"0000000011001111" when sig_inp <= "00101000011110101110" else
--"0000000011001011" when sig_inp <= "00101000101000111101" else
--"0000000011000111" when sig_inp <= "00101000110011001100" else
--"0000000011000011" when sig_inp <= "00101000111101011100" else
--"0000000010111111" when sig_inp <= "00101001000111101011" else
--"0000000010111100" when sig_inp <= "00101001010001111010" else
--"0000000010111000" when sig_inp <= "00101001011100001010" else
--"0000000010110100" when sig_inp <= "00101001100110011001" else
--"0000000010110001" when sig_inp <= "00101001110000101000" else
--"0000000010101101" when sig_inp <= "00101001111010111000" else
--"0000000010101010" when sig_inp <= "00101010000101000111" else
--"0000000010100110" when sig_inp <= "00101010001111010111" else
--"0000000010100011" when sig_inp <= "00101010011001100110" else
--"0000000010100000" when sig_inp <= "00101010100011110101" else
--"0000000010011101" when sig_inp <= "00101010101110000101" else
--"0000000010011010" when sig_inp <= "00101010111000010100" else
--"0000000010010110" when sig_inp <= "00101011000010100011" else
--"0000000010010011" when sig_inp <= "00101011001100110011" else
--"0000000010010001" when sig_inp <= "00101011010111000010" else
--"0000000010001110" when sig_inp <= "00101011100001010001" else
--"0000000010001011" when sig_inp <= "00101011101011100001" else
--"0000000010001000" when sig_inp <= "00101011110101110000" else
--"0000000010000101" when sig_inp <= "00101100000000000000" else
--"0000000010000011" when sig_inp <= "00101100001010001111" else
--"0000000010000000" when sig_inp <= "00101100010100011110" else
--"0000000001111110" when sig_inp <= "00101100011110101110" else
--"0000000001111011" when sig_inp <= "00101100101000111101" else
--"0000000001111001" when sig_inp <= "00101100110011001100" else
--"0000000001110110" when sig_inp <= "00101100111101011100" else
--"0000000001110100" when sig_inp <= "00101101000111101011" else
--"0000000001110010" when sig_inp <= "00101101010001111010" else
--"0000000001101111" when sig_inp <= "00101101011100001010" else
--"0000000001101101" when sig_inp <= "00101101100110011001" else
--"0000000001101011" when sig_inp <= "00101101110000101000" else
--"0000000001101001" when sig_inp <= "00101101111010111000" else
--"0000000001100111" when sig_inp <= "00101110000101000111" else
--"0000000001100101" when sig_inp <= "00101110001111010111" else
--"0000000001100011" when sig_inp <= "00101110011001100110" else
--"0000000001100001" when sig_inp <= "00101110100011110101" else
--"0000000001011111" when sig_inp <= "00101110101110000101" else
--"0000000001011101" when sig_inp <= "00101110111000010100" else
--"0000000001011011" when sig_inp <= "00101111000010100011" else
--"0000000001011001" when sig_inp <= "00101111001100110011" else
--"0000000001010111" when sig_inp <= "00101111010111000010" else
--"0000000001010110" when sig_inp <= "00101111100001010001" else
--"0000000001010100" when sig_inp <= "00101111101011100001" else
--"0000000001010010" when sig_inp <= "00101111110101110000" else
--"0000000001010001" when sig_inp <= "00110000000000000000" else
--"0000000001001111" when sig_inp <= "00110000001010001111" else
--"0000000001001110" when sig_inp <= "00110000010100011110" else
--"0000000001001100" when sig_inp <= "00110000011110101110" else
--"0000000001001010" when sig_inp <= "00110000101000111101" else
--"0000000001001001" when sig_inp <= "00110000110011001100" else
--"0000000001001000" when sig_inp <= "00110000111101011100" else
--"0000000001000110" when sig_inp <= "00110001000111101011" else
--"0000000001000101" when sig_inp <= "00110001010001111010" else
--"0000000001000011" when sig_inp <= "00110001011100001010" else
--"0000000001000010" when sig_inp <= "00110001100110011001" else
--"0000000001000001" when sig_inp <= "00110001110000101000" else
--"0000000000111111" when sig_inp <= "00110001111010111000" else
--"0000000000111110" when sig_inp <= "00110010000101000111" else
--"0000000000111101" when sig_inp <= "00110010001111010111" else
--"0000000000111100" when sig_inp <= "00110010011001100110" else
--"0000000000111010" when sig_inp <= "00110010100011110101" else
--"0000000000111001" when sig_inp <= "00110010101110000101" else
--"0000000000111000" when sig_inp <= "00110010111000010100" else
--"0000000000110111" when sig_inp <= "00110011000010100011" else
--"0000000000110110" when sig_inp <= "00110011001100110011" else
--"0000000000110101" when sig_inp <= "00110011010111000010" else
--"0000000000110100" when sig_inp <= "00110011100001010001" else
--"0000000000110011" when sig_inp <= "00110011101011100001" else
--"0000000000110010" when sig_inp <= "00110011110101110000" else
--"0000000000110001" when sig_inp <= "00110100000000000000" else
--"0000000000110000" when sig_inp <= "00110100001010001111" else
--"0000000000101111" when sig_inp <= "00110100010100011110" else
--"0000000000101110" when sig_inp <= "00110100011110101110" else
--"0000000000101101" when sig_inp <= "00110100101000111101" else
--"0000000000101100" when sig_inp <= "00110100110011001100" else
--"0000000000101011" when sig_inp <= "00110100111101011100" else
--"0000000000101010" when sig_inp <= "00110101000111101011" else
--"0000000000101001" when sig_inp <= "00110101010001111010" else
--"0000000000101001" when sig_inp <= "00110101011100001010" else
--"0000000000101000" when sig_inp <= "00110101100110011001" else
--"0000000000100111" when sig_inp <= "00110101110000101000" else
--"0000000000100110" when sig_inp <= "00110101111010111000" else
--"0000000000100101" when sig_inp <= "00110110000101000111" else
--"0000000000100101" when sig_inp <= "00110110001111010111" else
--"0000000000100100" when sig_inp <= "00110110011001100110" else
--"0000000000100011" when sig_inp <= "00110110100011110101" else
--"0000000000100011" when sig_inp <= "00110110101110000101" else
--"0000000000100010" when sig_inp <= "00110110111000010100" else
--"0000000000100001" when sig_inp <= "00110111000010100011" else
--"0000000000100001" when sig_inp <= "00110111001100110011" else
--"0000000000100000" when sig_inp <= "00110111010111000010" else
--"0000000000011111" when sig_inp <= "00110111100001010001" else
--"0000000000011111" when sig_inp <= "00110111101011100001" else
--"0000000000011110" when sig_inp <= "00110111110101110000" else
--"0000000000011101" when sig_inp <= "00111000000000000000" else
--"0000000000011101" when sig_inp <= "00111000001010001111" else
--"0000000000011100" when sig_inp <= "00111000010100011110" else
--"0000000000011100" when sig_inp <= "00111000011110101110" else
--"0000000000011011" when sig_inp <= "00111000101000111101" else
--"0000000000011011" when sig_inp <= "00111000110011001100" else
--"0000000000011010" when sig_inp <= "00111000111101011100" else
--"0000000000011001" when sig_inp <= "00111001000111101011" else
--"0000000000011001" when sig_inp <= "00111001010001111010" else
--"0000000000011000" when sig_inp <= "00111001011100001010" else
--"0000000000011000" when sig_inp <= "00111001100110011001" else
--"0000000000010111" when sig_inp <= "00111001110000101000" else
--"0000000000010111" when sig_inp <= "00111001111010111000" else
--"0000000000010111" when sig_inp <= "00111010000101000111" else
--"0000000000010110" when sig_inp <= "00111010001111010111" else
--"0000000000010110" when sig_inp <= "00111010011001100110" else
--"0000000000010101" when sig_inp <= "00111010100011110101" else
--"0000000000010101" when sig_inp <= "00111010101110000101" else
--"0000000000010100" when sig_inp <= "00111010111000010100" else
--"0000000000010100" when sig_inp <= "00111011000010100011" else
--"0000000000010100" when sig_inp <= "00111011001100110011" else
--"0000000000010011" when sig_inp <= "00111011010111000010" else
--"0000000000010011" when sig_inp <= "00111011100001010001" else
--"0000000000010010" when sig_inp <= "00111011101011100001" else
--"0000000000010010" when sig_inp <= "00111011110101110000" else
--"0000000000010010" when sig_inp <= "00111100000000000000" else
--"0000000000010001" when sig_inp <= "00111100001010001111" else
--"0000000000010001" when sig_inp <= "00111100010100011110" else
--"0000000000010001" when sig_inp <= "00111100011110101110" else
--"0000000000010000" when sig_inp <= "00111100101000111101" else
--"0000000000010000" when sig_inp <= "00111100110011001100" else
--"0000000000010000" when sig_inp <= "00111100111101011100" else
--"0000000000001111" when sig_inp <= "00111101000111101011" else
--"0000000000001111" when sig_inp <= "00111101010001111010" else
--"0000000000001111" when sig_inp <= "00111101011100001010" else
--"0000000000001110" when sig_inp <= "00111101100110011001" else
--"0000000000001110" when sig_inp <= "00111101110000101000" else
--"0000000000001110" when sig_inp <= "00111101111010111000" else
--"0000000000001101" when sig_inp <= "00111110000101000111" else
--"0000000000001101" when sig_inp <= "00111110001111010111" else
--"0000000000001101" when sig_inp <= "00111110011001100110" else
--"0000000000001101" when sig_inp <= "00111110100011110101" else
--"0000000000001100" when sig_inp <= "00111110101110000101" else
--"0000000000001100" when sig_inp <= "00111110111000010100" else
--"0000000000001100" when sig_inp <= "00111111000010100011" else
--"0000000000001100" when sig_inp <= "00111111001100110011" else
--"0000000000001011" when sig_inp <= "00111111010111000010" else
--"0000000000001011" when sig_inp <= "00111111100001010001" else
--"0000000000001011" when sig_inp <= "00111111101011100001" else
--"0000000000001011" when sig_inp <= "00111111110101110000" else
--"0000000000001010" when sig_inp <= "01000000000000000000" else
--"0000000000001010" when sig_inp <= "01000000001010001111" else
--"0000000000001010" when sig_inp <= "01000000010100011110" else
--"0000000000001010" when sig_inp <= "01000000011110101110" else
--"0000000000001010" when sig_inp <= "01000000101000111101" else
--"0000000000001001" when sig_inp <= "01000000110011001100" else
--"0000000000001001" when sig_inp <= "01000000111101011100" else
--"0000000000001001" when sig_inp <= "01000001000111101011" else
--"0000000000001001" when sig_inp <= "01000001010001111010" else
--"0000000000001001" when sig_inp <= "01000001011100001010" else
--"0000000000001000" when sig_inp <= "01000001100110011001" else
--"0000000000001000" when sig_inp <= "01000001110000101000" else
--"0000000000001000" when sig_inp <= "01000001111010111000" else
--"0000000000001000" when sig_inp <= "01000010000101000111" else
--"0000000000001000" when sig_inp <= "01000010001111010111" else
--"0000000000001000" when sig_inp <= "01000010011001100110" else
--"0000000000000111" when sig_inp <= "01000010100011110101" else
--"0000000000000111" when sig_inp <= "01000010101110000101" else
--"0000000000000111" when sig_inp <= "01000010111000010100" else
--"0000000000000111" when sig_inp <= "01000011000010100011" else
--"0000000000000111" when sig_inp <= "01000011001100110011" else
--"0000000000000111" when sig_inp <= "01000011010111000010" else
--"0000000000000111" when sig_inp <= "01000011100001010001" else
--"0000000000000110" when sig_inp <= "01000011101011100001" else
--"0000000000000110" when sig_inp <= "01000011110101110000" else
--"0000000000000110" when sig_inp <= "01000100000000000000" else
--"0000000000000110" when sig_inp <= "01000100001010001111" else
--"0000000000000110" when sig_inp <= "01000100010100011110" else
--"0000000000000110" when sig_inp <= "01000100011110101110" else
--"0000000000000110" when sig_inp <= "01000100101000111101" else
--"0000000000000110" when sig_inp <= "01000100110011001100" else
--"0000000000000101" when sig_inp <= "01000100111101011100" else
--"0000000000000101" when sig_inp <= "01000101000111101011" else
--"0000000000000101" when sig_inp <= "01000101010001111010" else
--"0000000000000101" when sig_inp <= "01000101011100001010" else
--"0000000000000101" when sig_inp <= "01000101100110011001" else
--"0000000000000101" when sig_inp <= "01000101110000101000" else
--"0000000000000101" when sig_inp <= "01000101111010111000" else
--"0000000000000101" when sig_inp <= "01000110000101000111" else
--"0000000000000101" when sig_inp <= "01000110001111010111" else
--"0000000000000100" when sig_inp <= "01000110011001100110" else
--"0000000000000100" when sig_inp <= "01000110100011110101" else
--"0000000000000100" when sig_inp <= "01000110101110000101" else
--"0000000000000100" when sig_inp <= "01000110111000010100" else
--"0000000000000100" when sig_inp <= "01000111000010100011" else
--"0000000000000100" when sig_inp <= "01000111001100110011" else
--"0000000000000100" when sig_inp <= "01000111010111000010" else
--"0000000000000100" when sig_inp <= "01000111100001010001" else
--"0000000000000100" when sig_inp <= "01000111101011100001" else
--"0000000000000100" when sig_inp <= "01000111110101110000" else
--"0000000000000100" when sig_inp <= "01001000000000000000" else
--"0000000000000011" when sig_inp <= "01001000001010001111" else
--"0000000000000011" when sig_inp <= "01001000010100011110" else
--"0000000000000011" when sig_inp <= "01001000011110101110" else
--"0000000000000011" when sig_inp <= "01001000101000111101" else
--"0000000000000011" when sig_inp <= "01001000110011001100" else
--"0000000000000011" when sig_inp <= "01001000111101011100" else
--"0000000000000011" when sig_inp <= "01001001000111101011" else
--"0000000000000011" when sig_inp <= "01001001010001111010" else
--"0000000000000011" when sig_inp <= "01001001011100001010" else
--"0000000000000011" when sig_inp <= "01001001100110011001" else
--"0000000000000011" when sig_inp <= "01001001110000101000" else
--"0000000000000011" when sig_inp <= "01001001111010111000" else
--"0000000000000011" when sig_inp <= "01001010000101000111" else
--"0000000000000011" when sig_inp <= "01001010001111010111" else
--"0000000000000010" when sig_inp <= "01001010011001100110" else
--"0000000000000010" when sig_inp <= "01001010100011110101" else
--"0000000000000010" when sig_inp <= "01001010101110000101" else
--"0000000000000010" when sig_inp <= "01001010111000010100" else
--"0000000000000010" when sig_inp <= "01001011000010100011" else
--"0000000000000010" when sig_inp <= "01001011001100110011" else
--"0000000000000010" when sig_inp <= "01001011010111000010" else
--"0000000000000010" when sig_inp <= "01001011100001010001" else
--"0000000000000010" when sig_inp <= "01001011101011100001" else
--"0000000000000010" when sig_inp <= "01001011110101110000" else
--"0000000000000010" when sig_inp <= "01001100000000000000" else
--"0000000000000010" when sig_inp <= "01001100001010001111" else
--"0000000000000010" when sig_inp <= "01001100010100011110" else
--"0000000000000010" when sig_inp <= "01001100011110101110" else
--"0000000000000010" when sig_inp <= "01001100101000111101" else
--"0000000000000010" when sig_inp <= "01001100110011001100" else
--"0000000000000010" when sig_inp <= "01001100111101011100" else
--"0000000000000010" when sig_inp <= "01001101000111101011" else
--"0000000000000010" when sig_inp <= "01001101010001111010" else
--"0000000000000010" when sig_inp <= "01001101011100001010" else
--"0000000000000010" when sig_inp <= "01001101100110011001" else
--"0000000000000001" when sig_inp <= "01001101110000101000" else
--"0000000000000001" when sig_inp <= "01001101111010111000" else
--"0000000000000001" when sig_inp <= "01001110000101000111" else
--"0000000000000001" when sig_inp <= "01001110001111010111" else
--"0000000000000001" when sig_inp <= "01001110011001100110" else
--"0000000000000001" when sig_inp <= "01001110100011110101" else
--"0000000000000001" when sig_inp <= "01001110101110000101" else
--"0000000000000001" when sig_inp <= "01001110111000010100" else
--"0000000000000001" when sig_inp <= "01001111000010100011" else
--"0000000000000001" when sig_inp <= "01001111001100110011" else
--"0000000000000001" when sig_inp <= "01001111010111000010" else
--"0000000000000001" when sig_inp <= "01001111100001010001" else
--"0000000000000001" when sig_inp <= "01001111101011100001" else
--"0000000000000001" when sig_inp <= "01001111110101110000" else
--"0000000000000001" when sig_inp <= "01010000000000000000" else
--"0000000000000001" when sig_inp <= "01010000001010001111" else
--"0000000000000001" when sig_inp <= "01010000010100011110" else
--"0000000000000001" when sig_inp <= "01010000011110101110" else
--"0000000000000001" when sig_inp <= "01010000101000111101" else
--"0000000000000001" when sig_inp <= "01010000110011001100" else
--"0000000000000001" when sig_inp <= "01010000111101011100" else
--"0000000000000001" when sig_inp <= "01010001000111101011" else
--"0000000000000001" when sig_inp <= "01010001010001111010" else
--"0000000000000001" when sig_inp <= "01010001011100001010" else
--"0000000000000001" when sig_inp <= "01010001100110011001" else
--"0000000000000001" when sig_inp <= "01010001110000101000" else
--"0000000000000000";

end Behavioral;
----------------------------------------------------------------------------------
